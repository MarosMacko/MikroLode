library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity UART_top is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity UART_top;

architecture RTL of UART_top is
	
begin

end architecture RTL;
