library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;

entity VGA_ROM is
    Port(clk, re     : in  STD_LOGIC;
         addr_tile   : in  STD_LOGIC_VECTOR(11 downto 0);
         addr_ship   : in  STD_LOGIC_VECTOR(12 downto 0);
         addr_hud    : in  STD_LOGIC_VECTOR(14 downto 0);
         output_hud  : out STD_LOGIC_VECTOR(3 downto 0);
         output_tile : out STD_LOGIC_VECTOR(3 downto 0);
         output_ship : out STD_LOGIC_VECTOR(3 downto 0));
end VGA_ROM;

architecture ROM of VGA_ROM is

    type Tile_ship_Rom_t is array (0 to 5887) of unsigned(3 downto 0);
    type Tile_tile_Rom_t is array (0 to 3327) of unsigned(3 downto 0);
    type HudRom_t is array (0 to 32767) of unsigned(3 downto 0);

    constant tile_ship_rom : Tile_ship_Rom_t := (
        x"3", x"3", x"C", x"C", x"C", x"C", x"F", x"E", x"E", x"C", x"C", x"C", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"F", x"E", x"E", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"C", x"E", x"E", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5",
        x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"C", x"C", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5",
        x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"3", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"3",
        x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"C", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"C", x"C", x"C", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5",
        x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"C", x"E", x"E", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"3", x"3", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3",
        x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"F", x"C", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"C", x"E", x"E", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"C", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"C", x"E", x"E", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"3", x"3", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"4", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5",
        x"3", x"3", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"3", x"3", x"3", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"8", x"4", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"3", x"3", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"3", x"3", x"B", x"E", x"E", x"C", x"C", x"C", x"C", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"3", x"3", x"B", x"E", x"E", x"C", x"E", x"C", x"C", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"3", x"3", x"B", x"E", x"E", x"C", x"E", x"C", x"E", x"C", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"3", x"3", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"5", x"3", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"3", x"3", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"3", x"3",
        x"3", x"3", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"3", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"8", x"4", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"B", x"8", x"8", x"8", x"8", x"A", x"C", x"9", x"8", x"8", x"4", x"B", x"E", x"E", x"E", x"B", x"8", x"8", x"8", x"8", x"B", x"B", x"9", x"8", x"8", x"3", x"3", x"B", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"B", x"E", x"E", x"A", x"8", x"8", x"8", x"4", x"B", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"B", x"E", x"E", x"E", x"A", x"9", x"3", x"3", x"B", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"B", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"B", x"8", x"8", x"8", x"8", x"A", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"8", x"8", x"9", x"D", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"B", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"9", x"B", x"E", x"E", x"E", x"E",
        x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"C", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"8", x"8", x"D", x"E", x"B", x"8", x"9", x"E", x"9", x"8", x"D", x"D", x"E", x"E", x"E", x"E", x"A", x"8", x"A", x"E", x"9", x"8", x"B", x"E", x"9", x"8", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"8", x"8", x"A", x"8", x"9", x"E", x"E", x"9", x"8", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"B", x"E", x"E", x"9", x"8", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"C", x"8", x"8", x"8", x"E", x"E", x"E", x"9", x"8", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"8", x"8", x"B", x"E", x"E", x"9", x"8", x"D", x"D",
        x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"8", x"A", x"E", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"8", x"8", x"E", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"9", x"8", x"A", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"A", x"8", x"9", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"A", x"A", x"8", x"B", x"9", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"A", x"D", x"8", x"9", x"9",
        x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"8", x"3", x"3", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"D", x"A", x"8", x"A", x"E", x"E", x"9", x"8", x"B", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"D", x"D", x"8", x"8", x"D", x"B", x"8", x"9", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"D", x"E", x"A", x"8", x"A", x"9", x"8", x"B", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"D", x"E", x"D", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"D", x"E", x"E", x"9", x"8", x"8", x"A", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"D", x"E", x"C", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5",
        x"8", x"4", x"B", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"D", x"E", x"E", x"E", x"A", x"9", x"3", x"3", x"B", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"B", x"E", x"E", x"9", x"8", x"8", x"8", x"4", x"B", x"E", x"E", x"E", x"B", x"8", x"8", x"8", x"8", x"A", x"A", x"9", x"8", x"8", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"B", x"8", x"8", x"8", x"8", x"B", x"D", x"A", x"8", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"D", x"9", x"8", x"8", x"A", x"E", x"E", x"9", x"8", x"8", x"8", x"4", x"B", x"E", x"E", x"E", x"9", x"8", x"B", x"D", x"9", x"B", x"E", x"9", x"8", x"D", x"3", x"3", x"B", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"D", x"8", x"4", x"B", x"E", x"E", x"E", x"9", x"8", x"9", x"A", x"E", x"E", x"E", x"9", x"8", x"D", x"3", x"3", x"B", x"E", x"E", x"E", x"C", x"9", x"8", x"8", x"9", x"D", x"E", x"9", x"8", x"D", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"B", x"9", x"8", x"9", x"E", x"9", x"8", x"8", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"B", x"8", x"9", x"E", x"9", x"8", x"D", x"8", x"4", x"B", x"E", x"E", x"B", x"9", x"B", x"E", x"A", x"8", x"A", x"E", x"9", x"8", x"D", x"3", x"3", x"B", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"A", x"E", x"E", x"9", x"8", x"D",
        x"C", x"E", x"E", x"E", x"B", x"8", x"9", x"B", x"8", x"9", x"E", x"E", x"9", x"8", x"D", x"D", x"9", x"D", x"E", x"E", x"9", x"8", x"B", x"E", x"9", x"8", x"A", x"E", x"9", x"8", x"D", x"D", x"8", x"9", x"C", x"B", x"8", x"9", x"E", x"E", x"B", x"8", x"8", x"E", x"9", x"8", x"D", x"D", x"8", x"8", x"A", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"B", x"E", x"E", x"A", x"8", x"8", x"B", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"C", x"8", x"8", x"D", x"E", x"9", x"8", x"8", x"9", x"E", x"E", x"E", x"8", x"8", x"D", x"E", x"E", x"9", x"8", x"B", x"D", x"8", x"9", x"9", x"8", x"E", x"E", x"E", x"8", x"8", x"D", x"E", x"E", x"9", x"8", x"B", x"A", x"8", x"B", x"A", x"8", x"A", x"E", x"E", x"8", x"8", x"D", x"D", x"C", x"8", x"8", x"E", x"9", x"8", x"E", x"B", x"8", x"9", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"9", x"C", x"D", x"8", x"9", x"E", x"E", x"8", x"8", x"E", x"E", x"8", x"8", x"D", x"A", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"8", x"8", x"A", x"E", x"8", x"8", x"D", x"E", x"E", x"E", x"E", x"9", x"8", x"C", x"E", x"E", x"B", x"8", x"9", x"E", x"8", x"8", x"D", x"E", x"E", x"E", x"C", x"8", x"9", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"8", x"8", x"D", x"E",
        x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"A", x"E", x"A", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"D", x"8", x"9", x"E", x"A", x"8", x"A", x"E", x"D", x"8", x"8", x"8", x"8", x"8", x"8", x"9", x"D", x"8", x"9", x"E", x"A", x"8", x"A", x"E", x"E", x"A", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"A", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"A", x"8", x"8", x"B", x"E", x"9", x"8", x"B", x"E", x"E", x"A", x"8", x"A", x"E", x"E", x"E", x"9", x"8", x"8", x"9", x"E", x"A", x"8", x"B", x"E", x"E", x"A", x"8", x"A", x"E", x"E", x"D", x"8", x"9", x"9", x"8", x"E", x"9", x"8", x"D", x"E", x"E", x"A", x"8", x"A", x"E", x"E", x"A", x"8", x"B", x"A", x"8", x"A", x"8", x"B", x"E", x"E", x"E", x"A", x"8", x"A", x"E", x"E", x"9", x"8", x"E", x"B", x"8", x"9", x"8", x"A", x"E", x"E", x"E", x"A", x"8", x"A", x"E", x"D", x"8", x"9", x"E", x"E", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"A", x"8", x"A", x"E", x"A", x"8", x"8", x"8", x"8", x"8", x"8", x"9", x"8", x"A", x"E", x"E", x"A", x"8", x"A", x"E", x"9", x"8", x"C", x"E", x"E", x"B", x"8", x"B", x"8", x"9", x"E", x"E", x"A", x"8", x"A", x"C", x"8", x"9", x"E", x"E", x"E", x"E", x"8",
        x"8", x"D", x"E", x"9", x"8", x"B", x"9", x"8", x"B", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"D", x"B", x"8", x"9", x"E", x"B", x"8", x"8", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"8", x"E", x"9", x"8", x"B", x"E", x"E", x"9", x"8", x"A", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"8", x"8", x"9", x"E", x"E", x"B", x"8", x"A", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"8", x"8", x"8", x"A", x"E", x"B", x"8", x"A", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"8", x"8", x"8", x"8", x"E", x"B", x"8", x"A", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"8", x"8", x"A", x"8", x"B", x"B", x"8", x"A", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"8", x"8", x"D", x"8", x"9", x"B", x"8", x"A", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"8", x"8", x"E", x"A", x"8", x"A", x"8", x"A", x"E", x"E", x"E", x"F", x"3", x"3", x"A", x"E", x"8", x"8", x"E", x"D", x"8", x"8", x"8", x"A", x"E", x"E", x"E", x"F", x"4", x"5", x"9", x"E", x"8", x"8", x"E", x"E", x"A", x"8", x"8", x"A", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"E", x"8", x"8", x"E", x"E", x"D", x"8", x"8", x"A", x"E", x"E", x"E", x"F", x"4", x"5",
        x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"B", x"8", x"E", x"E", x"E", x"8", x"A", x"E", x"E", x"9", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"B", x"8", x"E", x"9", x"A", x"E", x"E", x"9", x"9", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"8", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"A", x"E", x"E", x"B", x"9", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"8", x"B", x"8", x"E", x"E", x"E", x"8", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"9", x"9", x"E", x"B", x"8", x"E", x"E", x"9", x"9", x"3", x"3", x"B", x"E", x"E", x"E", x"9", x"9", x"E", x"E", x"E", x"9", x"9", x"E", x"E", x"9", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"9", x"E", x"E", x"9", x"8",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"E", x"E", x"9", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"E", x"8", x"E", x"E", x"8", x"E", x"E", x"8", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"8", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"A", x"E", x"E", x"E", x"E", x"9", x"A", x"E", x"E", x"E", x"E", x"E", x"9", x"E", x"E", x"A", x"8", x"B", x"8", x"E", x"E", x"9", x"A", x"B", x"8", x"E", x"E", x"E", x"9", x"8", x"8", x"8", x"E", x"E", x"9", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"E", x"E", x"A", x"8", x"8", x"9", x"E", x"E", x"9", x"8", x"8", x"9", x"E", x"E",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"B", x"B", x"8", x"E", x"E", x"9", x"A", x"E", x"8", x"E", x"E", x"8", x"B", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"A", x"B", x"9", x"E", x"E", x"9", x"A", x"B", x"9", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"E", x"B", x"9", x"E", x"E", x"9", x"9", x"B", x"9", x"E", x"A", x"E", x"E", x"9", x"9", x"E", x"E", x"B", x"9", x"E", x"E", x"9", x"A", x"B", x"9", x"E", x"A", x"E", x"8", x"A", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"8", x"B", x"E", x"8", x"E", x"E", x"A", x"8", x"8", x"8", x"8", x"A", x"E", x"A", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"8", x"8", x"8", x"B", x"E", x"A", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"8", x"B",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"8", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"9", x"A", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"9", x"A", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"8", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5",
        x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"8", x"B", x"E", x"8", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"8", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"9", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"A", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"B", x"8", x"E", x"E", x"E", x"9", x"A", x"B", x"8", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"A", x"8", x"8", x"8", x"9", x"E", x"E", x"9", x"8", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"4", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"3", x"3", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3",
        x"E", x"8", x"E", x"E", x"8", x"E", x"E", x"9", x"B", x"E", x"8", x"E", x"E", x"8", x"E", x"E", x"E", x"8", x"E", x"A", x"9", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"8", x"9", x"E", x"A", x"8", x"E", x"E", x"9", x"A", x"E", x"E", x"9", x"8", x"9", x"E", x"E", x"E", x"9", x"A", x"A", x"9", x"E", x"E", x"9", x"9", x"E", x"E", x"E", x"E", x"9", x"A", x"E", x"E", x"9", x"A", x"E", x"8", x"E", x"E", x"8", x"A", x"B", x"8", x"E", x"E", x"9", x"A", x"B", x"8", x"9", x"E", x"E", x"A", x"8", x"8", x"9", x"E", x"E", x"9", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3",
        x"9", x"A", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"8", x"B", x"E", x"E", x"8", x"8", x"B", x"8", x"8", x"8", x"9", x"E", x"B", x"9", x"E", x"E", x"9", x"A", x"E", x"9", x"E", x"8", x"B", x"8", x"E", x"E", x"9", x"A", x"B", x"9", x"E", x"E", x"9", x"9", x"E", x"E", x"E", x"8", x"B", x"E", x"E", x"E", x"9", x"9", x"B", x"9", x"E", x"E", x"9", x"A", x"E", x"E", x"E", x"8", x"B", x"8", x"E", x"E", x"8", x"B", x"E", x"8", x"E", x"E", x"8", x"B", x"E", x"E", x"E", x"8", x"B", x"9", x"8", x"8", x"9", x"E", x"E", x"A", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"8", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5",
        x"E", x"E", x"E", x"A", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"8", x"A", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"8", x"B", x"A", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"B", x"8", x"8", x"8", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"A", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"A", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"4", x"5", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"5", x"3", x"4", x"3", x"4", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"4", x"3", x"3", x"3", x"3", x"5", x"3", x"5", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"5", x"3", x"3", x"3",
        others => (others => '0'));
    constant tile_tile_rom : Tile_tile_Rom_t := (
        x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"2", x"2", x"8", x"E", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"2", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"A", x"3", x"3", x"3", x"3", x"A", x"3", x"3", x"3", x"3", x"A", x"3", x"3", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"C", x"7", x"6", x"3", x"3", x"C", x"7", x"6", x"3", x"3", x"C", x"7", x"6", x"3", x"3", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"3", x"1", x"1", x"0", x"F", x"3", x"1", x"1", x"0", x"F", x"3", x"1", x"1", x"0", x"F", x"3", x"3", x"2", x"2", x"3", x"F", x"3", x"2", x"2", x"3", x"F", x"3", x"2", x"2", x"3", x"F", x"3", x"3", x"4", x"4", x"5", x"F", x"3", x"4", x"4", x"5", x"F", x"3", x"4", x"4", x"5", x"F", x"3", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"7", x"7", x"6", x"F", x"3", x"3", x"3", x"B", x"F", x"F", x"3", x"3", x"B", x"F", x"F", x"3", x"3", x"B", x"F", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"B", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"3", x"3", x"3", x"3", x"F", x"3", x"3", x"3", x"3", x"F", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"3", x"3", x"3", x"F", x"6", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"1", x"0", x"F", x"F", x"3", x"7", x"6", x"F", x"F", x"8", x"E", x"3", x"3", x"3", x"2", x"B", x"1", x"0", x"F", x"F", x"B", x"7", x"6", x"F", x"F", x"A", x"F", x"2", x"3", x"3", x"2", x"3", x"1", x"0", x"F", x"F", x"3", x"7", x"6", x"F", x"F", x"3", x"3", x"2", x"3", x"3", x"2", x"B", x"1", x"0", x"F", x"F", x"B", x"7", x"6", x"F", x"F", x"3", x"3", x"2", x"3", x"3", x"2", x"3", x"1", x"0", x"F", x"F", x"3", x"7", x"6", x"F", x"F", x"8", x"E", x"2", x"3", x"3", x"2", x"3", x"3", x"0", x"F", x"F", x"3", x"F", x"6", x"F", x"F", x"A", x"F", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"F", x"F", x"3", x"3", x"3", x"F", x"F", x"3", x"3", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"3", x"8", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"3", x"3", x"2", x"3", x"3", x"2", x"A", x"A", x"4", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"A", x"A", x"2", x"3", x"3", x"2", x"2", x"F", x"5", x"5", x"5", x"0", x"7", x"5", x"5", x"5", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"8", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"3", x"3", x"3", x"3", x"3", x"A", x"A", x"A", x"4", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"A", x"A", x"A", x"3", x"3", x"3", x"F", x"F", x"5", x"5", x"5", x"0", x"7", x"5", x"5", x"5", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"8", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"3", x"3", x"3", x"3", x"3", x"A", x"A", x"A", x"4", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"A", x"A", x"A", x"3", x"3", x"3", x"F", x"F", x"5", x"5", x"5", x"0", x"7", x"5", x"5", x"5", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"8", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"3", x"3", x"3", x"3", x"3", x"A", x"A", x"A", x"4", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"A", x"A", x"A", x"3", x"3", x"3", x"F", x"F", x"5", x"5", x"5", x"0", x"7", x"5", x"5", x"5", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"C", x"7", x"7", x"1", x"2", x"4", x"7", x"7", x"3", x"3", x"3", x"3", x"3", x"A", x"A", x"A", x"7", x"7", x"7", x"1", x"2", x"4", x"7", x"7", x"A", x"A", x"A", x"3", x"3", x"3", x"F", x"F", x"6", x"6", x"6", x"0", x"3", x"5", x"6", x"6", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"8", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"3", x"3", x"3", x"3", x"3", x"A", x"A", x"A", x"4", x"4", x"4", x"1", x"5", x"4", x"4", x"4", x"A", x"A", x"A", x"3", x"3", x"3", x"F", x"F", x"5", x"5", x"5", x"0", x"7", x"5", x"5", x"5", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"C", x"1", x"1", x"7", x"2", x"4", x"1", x"1", x"3", x"3", x"3", x"3", x"3", x"A", x"A", x"A", x"1", x"1", x"1", x"7", x"2", x"4", x"1", x"1", x"A", x"A", x"A", x"3", x"3", x"3", x"F", x"F", x"0", x"0", x"0", x"6", x"3", x"5", x"0", x"0", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"1", x"1", x"1", x"3", x"3", x"3", x"3", x"3", x"4", x"4", x"4", x"3", x"3", x"3", x"3", x"1", x"C", x"C", x"C", x"1", x"3", x"3", x"2", x"2", x"5", x"5", x"5", x"3", x"3", x"3", x"1", x"C", x"B", x"C", x"C", x"C", x"1", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"1", x"C", x"C", x"C", x"C", x"C", x"1", x"3", x"2", x"3", x"7", x"7", x"7", x"2", x"3", x"3", x"1", x"C", x"C", x"C", x"C", x"C", x"1", x"F", x"2", x"2", x"6", x"6", x"6", x"3", x"3", x"3", x"3", x"1", x"C", x"C", x"C", x"1", x"F", x"F", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"1", x"1", x"1", x"F", x"F", x"3", x"2", x"B", x"B", x"B", x"E", x"2", x"3", x"3", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"B", x"C", x"C", x"F", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"B", x"C", x"B", x"F", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"B", x"C", x"C", x"F", x"3", x"3", x"3", x"2", x"8", x"E", x"2", x"2", x"2", x"8", x"E", x"3", x"B", x"C", x"B", x"F", x"3", x"3", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"A", x"F", x"3", x"B", x"C", x"C", x"F", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"E", x"F", x"F", x"F", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"8", x"E", x"2", x"8", x"E", x"2", x"3", x"3", x"2", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"F", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"F", x"3", x"3", x"3", x"2", x"3", x"3", x"7", x"7", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"3", x"3", x"3", x"A", x"B", x"B", x"5", x"5", x"6", x"5", x"5", x"5", x"5", x"5", x"5", x"7", x"F", x"F", x"3", x"B", x"F", x"F", x"7", x"7", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"3", x"2", x"3", x"3", x"7", x"7", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"3", x"A", x"B", x"B", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"F", x"F", x"3", x"B", x"F", x"F", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"F", x"F", x"3", x"2", x"2", x"3", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"F", x"F", x"3", x"2", x"2", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3",
        x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"E", x"F", x"3", x"F", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"3", x"3", x"3", x"3", x"2", x"8", x"A", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"E", x"F", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"8", x"A", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"2", x"2", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"3", x"2", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"3", x"2", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"3", x"2", x"3", x"0", x"1", x"9", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"3", x"2", x"3", x"F", x"1", x"1", x"1", x"1", x"0", x"0", x"0", x"F", x"F", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"3", x"B", x"F", x"F", x"B", x"F", x"F", x"F", x"F", x"3", x"3", x"2", x"3", x"3", x"2", x"3", x"3", x"B", x"F", x"3", x"B", x"F", x"F", x"F", x"F", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"B", x"2", x"A", x"B", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3",
        x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"0", x"0", x"2", x"8", x"E", x"2", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"0", x"8", x"9", x"0", x"A", x"F", x"2", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"1", x"8", x"0", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"3", x"3", x"0", x"8", x"9", x"0", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"2", x"3", x"3", x"3", x"3", x"0", x"9", x"1", x"0", x"2", x"2", x"3", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"3", x"2", x"1", x"8", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"2", x"0", x"1", x"8", x"1", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"0", x"1", x"A", x"8", x"1", x"8", x"0", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"0", x"1", x"A", x"8", x"1", x"0", x"3", x"0", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"2", x"1", x"8", x"1", x"0", x"0", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"2", x"2", x"8", x"0", x"0", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"2", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3",
        x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"2", x"0", x"0", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"0", x"8", x"0", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"2", x"3", x"0", x"9", x"8", x"0", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"3", x"2", x"0", x"1", x"8", x"1", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"0", x"1", x"1", x"0", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"0", x"8", x"0", x"2", x"2", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"0", x"9", x"9", x"0", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"2", x"0", x"9", x"0", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"2", x"2", x"8", x"E", x"0", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"2", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3",
        x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"2", x"2", x"0", x"0", x"1", x"1", x"2", x"0", x"1", x"0", x"E", x"2", x"3", x"3", x"2", x"2", x"3", x"0", x"1", x"9", x"8", x"8", x"1", x"A", x"9", x"0", x"F", x"2", x"3", x"3", x"2", x"3", x"0", x"A", x"8", x"A", x"0", x"1", x"8", x"8", x"0", x"2", x"2", x"2", x"3", x"3", x"2", x"0", x"1", x"8", x"0", x"0", x"3", x"0", x"0", x"0", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"0", x"1", x"8", x"0", x"0", x"0", x"1", x"0", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"0", x"1", x"8", x"8", x"1", x"9", x"8", x"1", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"0", x"1", x"8", x"8", x"A", x"1", x"8", x"1", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"0", x"1", x"8", x"0", x"0", x"2", x"1", x"8", x"0", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"0", x"A", x"A", x"0", x"3", x"3", x"3", x"0", x"3", x"2", x"2", x"3", x"3", x"3", x"2", x"2", x"1", x"8", x"1", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"2", x"2", x"8", x"0", x"0", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"2", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3",
        x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"0", x"E", x"2", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"1", x"0", x"2", x"3", x"3", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"0", x"1", x"8", x"8", x"1", x"2", x"3", x"3", x"2", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"0", x"8", x"8", x"1", x"0", x"2", x"3", x"3", x"2", x"3", x"2", x"3", x"3", x"3", x"0", x"0", x"9", x"8", x"1", x"0", x"2", x"3", x"3", x"3", x"2", x"3", x"2", x"2", x"0", x"0", x"0", x"A", x"8", x"1", x"0", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"0", x"0", x"1", x"8", x"8", x"8", x"1", x"0", x"2", x"3", x"3", x"3", x"3", x"2", x"2", x"0", x"1", x"9", x"8", x"9", x"1", x"9", x"9", x"1", x"0", x"2", x"3", x"3", x"3", x"3", x"0", x"1", x"8", x"8", x"1", x"0", x"0", x"0", x"1", x"8", x"8", x"0", x"3", x"3", x"3", x"2", x"0", x"9", x"9", x"0", x"0", x"3", x"3", x"3", x"0", x"0", x"9", x"1", x"2", x"3", x"2", x"2", x"8", x"0", x"0", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"0", x"0", x"2", x"2", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3",
        x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"8", x"E", x"2", x"3", x"3", x"2", x"2", x"3", x"0", x"0", x"3", x"3", x"3", x"0", x"0", x"1", x"1", x"0", x"2", x"3", x"3", x"2", x"3", x"0", x"A", x"1", x"0", x"0", x"0", x"1", x"8", x"8", x"9", x"0", x"2", x"3", x"3", x"2", x"3", x"0", x"1", x"8", x"8", x"1", x"1", x"8", x"8", x"1", x"0", x"2", x"2", x"3", x"3", x"2", x"3", x"0", x"1", x"8", x"9", x"8", x"8", x"8", x"0", x"0", x"2", x"2", x"3", x"3", x"3", x"2", x"0", x"1", x"8", x"1", x"0", x"0", x"8", x"9", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"8", x"1", x"0", x"2", x"1", x"8", x"1", x"0", x"2", x"2", x"3", x"3", x"3", x"3", x"0", x"1", x"8", x"0", x"3", x"3", x"1", x"8", x"1", x"1", x"0", x"2", x"2", x"3", x"3", x"3", x"0", x"1", x"8", x"0", x"3", x"3", x"0", x"9", x"8", x"8", x"8", x"0", x"2", x"3", x"3", x"3", x"2", x"0", x"8", x"1", x"3", x"3", x"3", x"0", x"0", x"0", x"8", x"1", x"2", x"2", x"3", x"2", x"2", x"8", x"0", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"0", x"0", x"E", x"2", x"2", x"3", x"2", x"A", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"A", x"F", x"2", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"2", x"3", x"3", x"3", x"2", x"2", x"2", x"2", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"2", x"2", x"3", x"3", x"3", x"3", x"2", x"3", x"3", x"3",
        others => (others => '0'));

    constant hud_rom : HudRom_t := (
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"7", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"F", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"A", x"C", x"C", x"C", x"C", x"C", x"C", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"4", x"4", x"4", x"4", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"7", x"7", x"7", x"4", x"4", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"7", x"7", x"7", x"7", x"4", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"7", x"7", x"7", x"4", x"4",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"C", x"C", x"C", x"C", x"C", x"C", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"4", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"4", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"0", x"0", x"0", x"4", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"0", x"0", x"0", x"4",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"C", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"9", x"A", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"4", x"4", x"4", x"0", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"4", x"0", x"4", x"0", x"0", x"4", x"4", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"4", x"0", x"0", x"0", x"0", x"0", x"4", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"4", x"0", x"0", x"0", x"0", x"4", x"4", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"E", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"E", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"8", x"7", x"6", x"9", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"8", x"7", x"6", x"9", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"3", x"3", x"1", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"3", x"3", x"1", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"5", x"5", x"7", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"4", x"4", x"5", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"4", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"4", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"4", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"4", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"4", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"4", x"4", x"4", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"D", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"D", x"D", x"4", x"F", x"D", x"D", x"4", x"4", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"D", x"D", x"4", x"4", x"F", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"F", x"4", x"4", x"F", x"F", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"F", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"D", x"D", x"F", x"4", x"F", x"4", x"4", x"F", x"D", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"D", x"D", x"4", x"4", x"4", x"F", x"F", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"4", x"D", x"4", x"4", x"4", x"F", x"F", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"4", x"4", x"F", x"D", x"D", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"D", x"D", x"4", x"D", x"F", x"F", x"F", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"4", x"4", x"D", x"D", x"D", x"D", x"8", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"4", x"4", x"4", x"D", x"D", x"D", x"9", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"4", x"D", x"D", x"D", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"4", x"4", x"4", x"4", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"D", x"F", x"F", x"4", x"4", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"D", x"D", x"4", x"4", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"4", x"4", x"4", x"4", x"F", x"F", x"D", x"D", x"D", x"D", x"B", x"B", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"7", x"2", x"2", x"2", x"F", x"2", x"2", x"7", x"7", x"7", x"7", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"2", x"2", x"2", x"F", x"2", x"2", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"8", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"B", x"B", x"D", x"D", x"8", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"8", x"9", x"D", x"D", x"9", x"B", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"D", x"D", x"8", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"D", x"D", x"9", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"D", x"B",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"F", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"B", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"F", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"B", x"D", x"B", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"F", x"D", x"B", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"E", x"F", x"D", x"B", x"D", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"B", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"E", x"F", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"E", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"D", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"F", x"D", x"B", x"B", x"B", x"D", x"B", x"D", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"F", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"F", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"B", x"D", x"B", x"D", x"B", x"D", x"D", x"D", x"B", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"6", x"6", x"D", x"D", x"D", x"6", x"6", x"D", x"D", x"D", x"D", x"6", x"6", x"6", x"D", x"D", x"6", x"6", x"F", x"D", x"D", x"6", x"6", x"F", x"0", x"0", x"6", x"6", x"F", x"F", x"D", x"D", x"6", x"6", x"F", x"D", x"D", x"6", x"6", x"F", x"0", x"0", x"6", x"F", x"F", x"0", x"D", x"D", x"7", x"7", x"F", x"D", x"D", x"7", x"7", x"F", x"0", x"0", x"7", x"7", x"0", x"0", x"D", x"D", x"7", x"7", x"F", x"0", x"0", x"7", x"7", x"F", x"0", x"0", x"0", x"7", x"7", x"7", x"D", x"D", x"5", x"5", x"F", x"0", x"0", x"5", x"5", x"F", x"0", x"0", x"0", x"0", x"5", x"5", x"D", x"D", x"5", x"5", x"F", x"0", x"0", x"5", x"5", x"F", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"4", x"4", x"F", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"4", x"0", x"0", x"D", x"D", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"0", x"4", x"4", x"4", x"D", x"D", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"0", x"F", x"0", x"0", x"F", x"F", x"F", x"D", x"D", x"4", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"4", x"4", x"4", x"F", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"4", x"4", x"F", x"F", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"6", x"0", x"0", x"0", x"6", x"0", x"0", x"0", x"0", x"6", x"0", x"0", x"0", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"F", x"0", x"0", x"0", x"6", x"F", x"0", x"0", x"6", x"F", x"0", x"0", x"F", x"F", x"0", x"6", x"F", x"0", x"0", x"0", x"6", x"F", x"0", x"0", x"6", x"F", x"0", x"0", x"0", x"0", x"0", x"7", x"F", x"0", x"0", x"0", x"7", x"F", x"0", x"0", x"7", x"F", x"0", x"0", x"0", x"0", x"0", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"0", x"0", x"7", x"F", x"0", x"5", x"5", x"F", x"F", x"5", x"F", x"F", x"F", x"F", x"5", x"F", x"0", x"0", x"5", x"F", x"0", x"5", x"5", x"F", x"D", x"5", x"F", x"0", x"0", x"0", x"5", x"F", x"0", x"0", x"5", x"F", x"0", x"4", x"4", x"F", x"D", x"4", x"F", x"0", x"0", x"0", x"4", x"F", x"0", x"F", x"4", x"F", x"D", x"4", x"F", x"F", x"0", x"4", x"F", x"0", x"0", x"0", x"4", x"F", x"F", x"F", x"4", x"F", x"D", x"F", x"F", x"0", x"0", x"0", x"F", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"F", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"2", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"7", x"7", x"7", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"F", x"7", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"7", x"7", x"7", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"6", x"6", x"6", x"6", x"6", x"D", x"D", x"D", x"D", x"6", x"6", x"6", x"6", x"D", x"D", x"D", x"6", x"F", x"F", x"F", x"6", x"6", x"D", x"D", x"6", x"6", x"F", x"F", x"6", x"6", x"D", x"D", x"6", x"F", x"0", x"0", x"0", x"6", x"F", x"D", x"6", x"F", x"F", x"D", x"D", x"F", x"F", x"D", x"7", x"F", x"0", x"0", x"0", x"7", x"F", x"0", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"F", x"0", x"0", x"7", x"7", x"F", x"0", x"0", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"5", x"5", x"5", x"5", x"5", x"F", x"F", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"D", x"D", x"5", x"F", x"F", x"F", x"F", x"F", x"0", x"0", x"0", x"0", x"0", x"F", x"5", x"5", x"F", x"D", x"4", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"0", x"0", x"4", x"4", x"F", x"D", x"4", x"F", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"F", x"F", x"D", x"D", x"F", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"F", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"F", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"F", x"B", x"B", x"B", x"B", x"B", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"0", x"0", x"0", x"0", x"0", x"F", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"4", x"4", x"4", x"4", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"7", x"7", x"4", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"D", x"A", x"9", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"C", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"7", x"7", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"4", x"7", x"7", x"7", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"7", x"7", x"7", x"7", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"4", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"C", x"C", x"C", x"C", x"C", x"C", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"0", x"0", x"0", x"0", x"4", x"4", x"0", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"4", x"4", x"0", x"0", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"4", x"0", x"0", x"0", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"A", x"D", x"0", x"0", x"0", x"0", x"0", x"E", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"A", x"D", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"C", x"C", x"C", x"C", x"C", x"C", x"A", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"8", x"7", x"7", x"6", x"E", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"8", x"D", x"B", x"E", x"E", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"8", x"8", x"9", x"E", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"8", x"9", x"E", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"7", x"7", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"7", x"7", x"7", x"7", x"2", x"2", x"F", x"7", x"7", x"7", x"7", x"2", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"2", x"2", x"2", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"8", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"E", x"F", x"D", x"D", x"9", x"B", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"9", x"B", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"B", x"E", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"B", x"B", x"D", x"E", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"D", x"E", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"E", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"2", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"F", x"F", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"F", x"2", x"2", x"F", x"F", x"F", x"2", x"F", x"F", x"F", x"2", x"2", x"2", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"2", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"F", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"2", x"2", x"F", x"F", x"2", x"2", x"2", x"2", x"F", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"2", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"F", x"F", x"F", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"2", x"2", x"2", x"F", x"F", x"F", x"2", x"2", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"8", x"8", x"8", x"8", x"8", x"8", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"8", x"8", x"8", x"8", x"8", x"D", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"D", x"9", x"D", x"9", x"9", x"8", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"D", x"8", x"D", x"B", x"9", x"9", x"9", x"B", x"8", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"8", x"B", x"9", x"9", x"9", x"E", x"E", x"D", x"8", x"D", x"D", x"D", x"D", x"D", x"D", x"B", x"8", x"B", x"9", x"9", x"9", x"E", x"E", x"D", x"8", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"9", x"9", x"9", x"E", x"E", x"E", x"D", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"8", x"9", x"9", x"E", x"E", x"E", x"E", x"D", x"9", x"D", x"D", x"D", x"B", x"B", x"B", x"D", x"8", x"9", x"9", x"E", x"E", x"E", x"E", x"D", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"B", x"8", x"9", x"E", x"E", x"E", x"E", x"E", x"D", x"9", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"8", x"D", x"E", x"E", x"E", x"E", x"D", x"9", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"8", x"D", x"9", x"E", x"D", x"D", x"9", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"8", x"D", x"9", x"E", x"D", x"D", x"9", x"D", x"D", x"D", x"D", x"B", x"D", x"D", x"D", x"D", x"8", x"9", x"9", x"9", x"9", x"9", x"B", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"F", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"B", x"B", x"B", x"B", x"B", x"0", x"0", x"0", x"0", x"0", x"F", x"B", x"B", x"B", x"B", x"B", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0",
        x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"B", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"0", x"0", x"0", x"0", x"F", x"F", x"F", x"B", x"0", x"0", x"0", x"F", x"F", x"F", x"F", x"0", x"0", x"0", x"0", x"F", x"F", x"B", x"B", x"D", x"D", x"F", x"F", x"F", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"0", x"0", x"0", x"0", x"0", x"0", x"F", x"F", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"F", x"0", x"0", x"F", x"F", x"F", x"D", x"D", x"D", x"0",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"9", x"F", x"9", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"9", x"9", x"9", x"F", x"F", x"9", x"F", x"F", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"8", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"8", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"A", x"9", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"8", x"A", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"A", x"9", x"9", x"9", x"9", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"9", x"9", x"9", x"9", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"A", x"9", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4",
        x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"8", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"F", x"F", x"8", x"8", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"5", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"F", x"F", x"F", x"5", x"5", x"4", x"4", x"4", x"4", x"4", x"F", x"4", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"5", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"5", x"F", x"F",
        x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"4", x"8", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"8", x"8", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"8", x"9", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"8", x"9", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"8", x"9", x"9", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"F", x"F", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"F", x"F", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F",
        x"8", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"9", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"9", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"8", x"8", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"8", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"8", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"8", x"8", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"8", x"8", x"8", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"8", x"8", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"5",
        x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"9", x"9", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"9", x"9", x"9", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"E", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"E", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"E", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"E", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"E", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"E", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"5", x"5",
        x"9", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"9", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"9", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"9", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"8", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E",
        x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E",
        x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"8", x"5", x"5", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"F", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"5", x"5", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"5", x"8", x"4", x"4", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"4", x"4", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"4", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"8", x"5", x"5", x"5", x"5", x"5", x"5", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"5", x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"5", x"5", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"5", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"5", x"5", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"8", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"F", x"F", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E", x"E", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"E", x"8", x"E", x"E", x"E",
        x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"E", x"8", x"E",
        x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"9", x"9", x"9", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"9", x"9", x"9", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D", x"D",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"7", x"7", x"7", x"7", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"F", x"4", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"4", x"4", x"4", x"4", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F", x"F",
        others => (others => '0'));

begin

    tile_ship_rom_process : process(clk)
    begin
        if (rising_edge(clk)) then
            if (re = '1') then
                output_ship <= std_logic_vector(tile_ship_rom(to_integer(unsigned(addr_ship))));
            end if;
        end if;
    end process;

    tile_tile_rom_process : process(clk)
    begin
        if (rising_edge(clk)) then
            if (re = '1') then
                output_tile <= std_logic_vector(tile_tile_rom(to_integer(unsigned(addr_tile))));
            end if;
        end if;
    end process;

    hud_rom_process : process(clk)
    begin
        if (rising_edge(clk)) then
            if (re = '1') then
                output_hud <= std_logic_vector(hud_rom(to_integer(unsigned(addr_hud))));
            end if;
        end if;
    end process;

end ROM;

