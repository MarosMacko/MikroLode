library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity VGA_pixel_gen is
    Port(clk         : in  STD_LOGIC;
         pixel_x     : in  STD_LOGIC_VECTOR(10 downto 0);
         pixel_y     : in  STD_LOGIC_VECTOR(10 downto 0);
         RAM_address : out STD_LOGIC_VECTOR(10 downto 0);
         RAM_data    : in  STD_LOGIC_VECTOR(8 downto 0);
         R, G, B     : out STD_LOGIC_VECTOR(6 downto 0));
end VGA_pixel_gen;

architecture Behavioral of VGA_pixel_gen is
    --signal R_int, G_int, B_int : STD_LOGIC_VECTOR(7 downto 0) := (others => '0');
    signal re : std_logic := '1';
    type RomType is array (0 to 4095) of unsigned(7 downto 0);

    constant r_rom : RomType := (
        X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7d", X"7d", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7e", X"7f", X"7e", X"79", X"5a", X"4e", X"78", X"7e", X"7f", X"7f", X"7f", X"7b", X"7e", X"7e", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7d", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7a", X"23", X"00", X"00", X"1c", X"78", X"7a", X"7f", X"7f", X"7f", X"7e", X"7a", X"7d", X"7e", X"7e", X"7e", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"78", X"12", X"00", X"00", X"00", X"00", X"02", X"5f", X"7a", X"7e", X"7f", X"7e", X"7e", X"7e", X"7e", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"69", X"00", X"00", X"01", X"00", X"00", X"02", X"00", X"00", X"2e", X"77", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"47", X"00", X"00", X"00", X"02", X"02", X"01", X"02", X"00", X"00", X"00", X"16", X"78", X"7d", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"76", X"25", X"00", X"00", X"00", X"02", X"00", X"00", X"00", X"02", X"01", X"00", X"00", X"00", X"00", X"79", X"7c", X"7f", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"79", X"12", X"00", X"01", X"01", X"03", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"01", X"00", X"02", X"01", X"59", X"77", X"7e", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"72", X"15", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"58", X"7e", X"7f", X"7d", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"79", X"05", X"00", X"00", X"00", X"01", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"04", X"4c", X"77", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"76", X"0a", X"01", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"01", X"00", X"00", X"00", X"00", X"03", X"01", X"00", X"40", X"7a", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7c", X"0a", X"00", X"00", X"00", X"02", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"50", X"78", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"74", X"09", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"02", X"00", X"4c", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"79", X"1c", X"00", X"00", X"01", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"66", X"7a", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"75", X"25", X"02", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"02", X"03", X"00", X"75", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"4c", X"00", X"00", X"00", X"00", X"01", X"02", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"01", X"05", X"02", X"00", X"00", X"08", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7e", X"7f", X"7d", X"7a", X"68", X"02", X"00", X"00", X"00", X"01", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"0d", X"19", X"27", X"2e", X"2c", X"23", X"17", X"0a", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"10", X"72", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7d", X"76", X"03", X"00", X"00", X"00", X"02", X"01", X"00", X"03", X"00", X"00", X"23", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7c", X"23", X"00", X"00", X"03", X"00", X"00", X"04", X"02", X"03", X"00", X"00", X"36", X"7c", X"7d", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"79", X"0f", X"01", X"02", X"01", X"03", X"01", X"02", X"00", X"05", X"61", X"7c", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"76", X"27", X"56", X"78", X"7f", X"7e", X"7f", X"7c", X"78", X"64", X"03", X"00", X"02", X"00", X"00", X"00", X"00", X"00", X"01", X"69", X"7a", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"79", X"3b", X"01", X"00", X"01", X"00", X"00", X"00", X"01", X"41", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"77", X"72", X"12", X"00", X"02", X"7a", X"7d", X"7f", X"7f", X"7f", X"7f", X"7c", X"78", X"41", X"00", X"00", X"03", X"00", X"00", X"02", X"00", X"08", X"78", X"7b", X"7f", X"7e", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7c", X"73", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"78", X"7c", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"0b", X"00", X"00", X"00", X"5a", X"77", X"7c", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7d", X"0b", X"00", X"00", X"00", X"00", X"02", X"00", X"14", X"7c", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7a", X"06", X"00", X"01", X"00", X"02", X"02", X"27", X"7a", X"7f", X"7f", X"7b", X"7e", X"7f", X"7f", X"7f", X"7b", X"77", X"0b", X"00", X"00", X"02", X"05", X"0a", X"75", X"7e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"77", X"29", X"00", X"00", X"01", X"00", X"01", X"00", X"6d", X"79", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"77", X"3a", X"00", X"00", X"00", X"00", X"00", X"0b", X"78", X"7d", X"7f", X"7f", X"7d", X"7a", X"7d", X"7d", X"7f", X"7b", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"4b", X"7c", X"7f", X"7f", X"7e", X"7e", X"7d", X"7f", X"7e", X"7f", X"7d", X"10", X"00", X"00", X"01", X"00", X"00", X"00", X"78", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"68", X"00", X"00", X"03", X"01", X"00", X"16", X"73", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"78", X"59", X"01", X"00", X"03", X"01", X"02", X"01", X"00", X"00", X"06", X"7a", X"7d", X"7d", X"7e", X"7f", X"7d", X"7f", X"7e", X"7e", X"7a", X"73", X"1a", X"00", X"00", X"00", X"00", X"00", X"36", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7e", X"79", X"0d", X"00", X"00", X"00", X"00", X"08", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7a", X"4f", X"01", X"00", X"01", X"05", X"02", X"01", X"00", X"02", X"01", X"01", X"65", X"78", X"7b", X"7c", X"7c", X"7d", X"7f", X"7f", X"7d", X"7e", X"7f", X"7c", X"06", X"00", X"01", X"02", X"01", X"03", X"7a", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7b", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7e", X"7f", X"7f", X"7c", X"76", X"3e", X"02", X"03", X"00", X"00", X"00", X"6f", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"78", X"37", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"02", X"00", X"04", X"03", X"08", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7e", X"7d", X"78", X"01", X"00", X"00", X"03", X"01", X"0c", X"78", X"7b", X"7d", X"7f", X"7f", X"7f", X"7e", X"7e", X"7c", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7a", X"7c", X"05", X"02", X"00", X"00", X"00", X"0f", X"76", X"7a", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"62", X"5b", X"62", X"61", X"1a", X"00", X"00", X"01", X"57", X"58", X"59", X"59", X"5e", X"77", X"7b", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"77", X"1a", X"03", X"00", X"00", X"00", X"01", X"76", X"7b", X"7f", X"7f", X"7f", X"7d", X"7d", X"7d", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"7f", X"7d", X"39", X"00", X"00", X"00", X"00", X"00", X"7c", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7b", X"09", X"00", X"00", X"45", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7a", X"7f", X"7f", X"7c", X"7c", X"04", X"00", X"00", X"00", X"00", X"23", X"7a", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7b", X"7c", X"7f", X"7f", X"7f", X"7c", X"02", X"00", X"01", X"00", X"00", X"1f", X"7c", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"75", X"30", X"00", X"01", X"06", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7b", X"7c", X"7f", X"7f", X"7f", X"7c", X"7c", X"7d", X"7f", X"7f", X"7f", X"7b", X"2f", X"00", X"00", X"01", X"00", X"00", X"78", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7b", X"7f", X"7f", X"7f", X"7d", X"7f", X"7c", X"73", X"27", X"00", X"00", X"02", X"01", X"00", X"67", X"7d", X"7f", X"7f", X"7f", X"7e", X"7c", X"7c", X"7c", X"7e", X"7f", X"7f", X"7d", X"64", X"00", X"00", X"00", X"05", X"77", X"7d", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"79", X"6a", X"00", X"01", X"00", X"00", X"00", X"1c", X"75", X"7c", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7b", X"79", X"78", X"04", X"01", X"00", X"01", X"02", X"03", X"79", X"7b", X"7c", X"7f", X"7f", X"7c", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7a", X"05", X"00", X"00", X"00", X"26", X"77", X"7d", X"7f", X"7f", X"7e", X"7c", X"7d", X"7f", X"7c", X"57", X"05", X"7d", X"7f", X"7f", X"7f", X"7f", X"7c", X"7d", X"7b", X"77", X"01", X"00", X"00", X"00", X"00", X"04", X"7b", X"7c", X"7f", X"7f", X"7d", X"7e", X"7b", X"7f", X"7f", X"7e", X"7b", X"7d", X"7a", X"3b", X"00", X"00", X"03", X"00", X"00", X"0d", X"77", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7c", X"78", X"19", X"00", X"00", X"00", X"02", X"76", X"7c", X"7d", X"7f", X"7f", X"7f", X"7d", X"76", X"23", X"03", X"00", X"02", X"78", X"7b", X"7b", X"7e", X"7f", X"7f", X"7f", X"7b", X"75", X"14", X"01", X"05", X"02", X"01", X"00", X"33", X"7c", X"7e", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7d", X"7b", X"02", X"01", X"00", X"00", X"00", X"02", X"59", X"7a", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7c", X"75", X"03", X"00", X"00", X"01", X"03", X"7f", X"7f", X"7f", X"7a", X"75", X"45", X"01", X"00", X"00", X"00", X"00", X"05", X"7f", X"7f", X"7f", X"7c", X"7d", X"7d", X"7f", X"7d", X"78", X"59", X"04", X"01", X"01", X"00", X"00", X"04", X"7b", X"7b", X"7c", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"77", X"57", X"00", X"00", X"01", X"00", X"04", X"06", X"77", X"7e", X"7d", X"7c", X"7b", X"7b", X"7e", X"7d", X"7f", X"7f", X"7f", X"7a", X"08", X"00", X"00", X"00", X"00", X"10", X"77", X"72", X"1c", X"00", X"00", X"04", X"01", X"00", X"00", X"00", X"01", X"01", X"7b", X"7b", X"7e", X"7f", X"7e", X"7f", X"7f", X"7d", X"7d", X"7a", X"00", X"01", X"00", X"01", X"02", X"01", X"60", X"7a", X"7c", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"78", X"14", X"00", X"01", X"01", X"00", X"00", X"00", X"7c", X"7f", X"7e", X"7f", X"7e", X"7e", X"7e", X"7e", X"7e", X"7b", X"74", X"4b", X"03", X"01", X"00", X"00", X"00", X"01", X"03", X"00", X"00", X"01", X"00", X"00", X"01", X"00", X"02", X"01", X"00", X"02", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7c", X"03", X"00", X"00", X"00", X"01", X"00", X"24", X"77", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7c", X"79", X"02", X"01", X"00", X"00", X"00", X"00", X"01", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7a", X"75", X"08", X"00", X"00", X"00", X"00", X"00", X"03", X"00", X"02", X"00", X"00", X"01", X"01", X"00", X"00", X"01", X"00", X"00", X"05", X"7b", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7a", X"07", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"79", X"28", X"00", X"00", X"00", X"00", X"00", X"02", X"07", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7b", X"36", X"00", X"00", X"02", X"05", X"03", X"02", X"00", X"04", X"00", X"00", X"00", X"07", X"01", X"00", X"03", X"00", X"02", X"00", X"0d", X"7b", X"7e", X"7d", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"07", X"00", X"00", X"00", X"00", X"00", X"00", X"46", X"7b", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7c", X"05", X"00", X"00", X"02", X"00", X"00", X"00", X"03", X"7d", X"7f", X"7e", X"7e", X"7e", X"7f", X"7d", X"7e", X"7f", X"7c", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"06", X"55", X"76", X"06", X"03", X"00", X"00", X"00", X"00", X"1a", X"77", X"7a", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7e", X"05", X"00", X"01", X"01", X"01", X"00", X"00", X"09", X"7d", X"7f", X"7e", X"7d", X"7d", X"7c", X"7d", X"7b", X"03", X"02", X"00", X"00", X"00", X"01", X"00", X"02", X"7a", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"75", X"41", X"02", X"00", X"04", X"00", X"02", X"00", X"00", X"00", X"00", X"45", X"7d", X"7d", X"7a", X"05", X"00", X"01", X"00", X"00", X"00", X"37", X"7b", X"7e", X"7f", X"7f", X"7e", X"7d", X"7d", X"7e", X"7f", X"7e", X"03", X"01", X"00", X"00", X"00", X"00", X"00", X"03", X"7b", X"7f", X"7f", X"7e", X"7f", X"7f", X"7b", X"4b", X"03", X"00", X"00", X"00", X"00", X"00", X"07", X"05", X"78", X"7a", X"7c", X"7d", X"7f", X"7f", X"7d", X"7b", X"7a", X"0a", X"02", X"00", X"00", X"00", X"00", X"01", X"03", X"52", X"7c", X"7e", X"7f", X"7b", X"4a", X"00", X"01", X"00", X"01", X"00", X"00", X"50", X"7b", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7d", X"7d", X"7c", X"02", X"01", X"00", X"00", X"00", X"00", X"00", X"02", X"75", X"7c", X"7d", X"7f", X"7f", X"7d", X"78", X"0d", X"03", X"04", X"00", X"00", X"00", X"00", X"02", X"01", X"45", X"78", X"7c", X"7f", X"7f", X"7f", X"7f", X"7d", X"43", X"00", X"00", X"00", X"00", X"00", X"10", X"4d", X"76", X"7e", X"7f", X"7f", X"7f", X"7a", X"14", X"00", X"00", X"02", X"01", X"02", X"03", X"77", X"7c", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"78", X"46", X"02", X"02", X"00", X"02", X"00", X"00", X"01", X"00", X"36", X"77", X"7c", X"7f", X"7b", X"7c", X"7b", X"04", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0b", X"78", X"7e", X"7f", X"7f", X"7d", X"7e", X"7b", X"0a", X"00", X"00", X"00", X"3c", X"78", X"7b", X"7f", X"7f", X"7f", X"7e", X"7c", X"7f", X"7a", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"79", X"7c", X"7d", X"7e", X"7d", X"7d", X"7f", X"7e", X"7c", X"77", X"0a", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"03", X"02", X"79", X"7c", X"7f", X"7f", X"7c", X"61", X"00", X"00", X"00", X"02", X"02", X"00", X"00", X"00", X"00", X"04", X"7a", X"7c", X"7f", X"7f", X"7f", X"7f", X"79", X"2b", X"53", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"75", X"0d", X"00", X"00", X"02", X"05", X"00", X"01", X"08", X"78", X"7c", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"79", X"77", X"03", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"02", X"77", X"7f", X"7f", X"7f", X"7b", X"35", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"03", X"00", X"5a", X"7d", X"7e", X"7e", X"7c", X"7e", X"7f", X"7f", X"7f", X"7d", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7c", X"7c", X"7a", X"03", X"02", X"06", X"00", X"00", X"00", X"00", X"0f", X"74", X"7c", X"7f", X"7d", X"7c", X"7e", X"7e", X"7d", X"7c", X"64", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"02", X"00", X"62", X"7d", X"7f", X"7e", X"7a", X"16", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"03", X"02", X"00", X"16", X"79", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"78", X"0c", X"00", X"00", X"00", X"02", X"01", X"06", X"00", X"22", X"76", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"1f", X"00", X"00", X"01", X"00", X"00", X"00", X"02", X"00", X"00", X"00", X"34", X"7e", X"7f", X"7f", X"7b", X"09", X"00", X"00", X"02", X"03", X"02", X"00", X"00", X"00", X"00", X"00", X"02", X"73", X"75", X"7d", X"7f", X"7e", X"7e", X"7d", X"7e", X"7b", X"7c", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"7c", X"5d", X"03", X"03", X"01", X"02", X"01", X"00", X"00", X"00", X"49", X"77", X"7c", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7a", X"00", X"00", X"00", X"00", X"03", X"00", X"01", X"03", X"00", X"00", X"00", X"1e", X"79", X"7f", X"7e", X"7b", X"04", X"00", X"00", X"00", X"00", X"01", X"01", X"00", X"00", X"00", X"00", X"00", X"0b", X"77", X"7b", X"7c", X"7c", X"7d", X"7f", X"7f", X"7f", X"7e", X"7e", X"7b", X"7f", X"7f", X"7f", X"7c", X"78", X"07", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"76", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7c", X"7a", X"0e", X"00", X"00", X"01", X"00", X"00", X"00", X"02", X"00", X"00", X"00", X"00", X"0c", X"7c", X"7f", X"7f", X"7c", X"01", X"00", X"00", X"02", X"03", X"01", X"00", X"00", X"00", X"01", X"01", X"02", X"00", X"4c", X"7b", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7c", X"7d", X"79", X"1b", X"00", X"00", X"00", X"02", X"03", X"00", X"00", X"00", X"07", X"7c", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7b", X"5e", X"00", X"01", X"01", X"00", X"00", X"00", X"00", X"02", X"01", X"00", X"00", X"00", X"06", X"7b", X"7c", X"78", X"6d", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"79", X"7e", X"7d", X"7e", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"79", X"60", X"00", X"00", X"01", X"00", X"00", X"02", X"00", X"00", X"00", X"2f", X"79", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"03", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"7e", X"7f", X"76", X"3e", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"75", X"7e", X"7f", X"7c", X"7f", X"7f", X"7e", X"7f", X"7f", X"7c", X"7c", X"79", X"04", X"02", X"00", X"00", X"00", X"03", X"01", X"00", X"01", X"03", X"7a", X"7d", X"7e", X"7c", X"7a", X"7e", X"7c", X"77", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"01", X"00", X"03", X"00", X"00", X"00", X"03", X"79", X"7c", X"72", X"27", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0b", X"7c", X"7f", X"7f", X"7c", X"7b", X"7b", X"7c", X"7f", X"7f", X"7b", X"08", X"00", X"00", X"01", X"02", X"03", X"00", X"00", X"01", X"00", X"03", X"7b", X"7f", X"7f", X"7d", X"7f", X"7f", X"7c", X"0a", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"00", X"58", X"77", X"72", X"13", X"00", X"01", X"02", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"05", X"00", X"08", X"75", X"7d", X"7f", X"7e", X"7f", X"7f", X"7b", X"77", X"0d", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"03", X"26", X"76", X"7c", X"7f", X"7f", X"7c", X"78", X"0c", X"00", X"01", X"00", X"00", X"00", X"00", X"01", X"01", X"00", X"00", X"00", X"01", X"01", X"00", X"00", X"00", X"36", X"72", X"72", X"07", X"00", X"00", X"01", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"01", X"00", X"06", X"68", X"7b", X"7d", X"7f", X"7f", X"7c", X"11", X"00", X"00", X"01", X"00", X"02", X"03", X"01", X"00", X"00", X"00", X"03", X"7f", X"7f", X"7d", X"7a", X"79", X"65", X"06", X"00", X"02", X"03", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"00", X"00", X"00", X"00", X"18", X"71", X"79", X"04", X"04", X"00", X"00", X"00", X"00", X"02", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"2b", X"7b", X"7d", X"78", X"08", X"02", X"00", X"03", X"04", X"01", X"00", X"00", X"00", X"01", X"00", X"00", X"2a", X"7a", X"7e", X"7f", X"7d", X"2d", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"01", X"00", X"00", X"0a", X"75", X"7e", X"7b", X"12", X"00", X"00", X"00", X"00", X"01", X"02", X"02", X"00", X"00", X"00", X"00", X"00", X"01", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"26", X"72", X"3e", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"01", X"00", X"00", X"00", X"73", X"7a", X"79", X"26", X"00", X"00", X"04", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0d", X"7a", X"7c", X"7f", X"7f", X"78", X"6f", X"0b", X"00", X"00", X"01", X"03", X"03", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"04", X"04", X"03", X"00", X"00", X"0e", X"23", X"1b", X"1d", X"02", X"00", X"01", X"01", X"00", X"00", X"00", X"03", X"3a", X"15", X"00", X"00", X"00", X"00", X"00", X"00", X"02", X"01", X"03", X"01", X"00", X"00", X"00", X"00", X"00", X"01", X"01", X"01", X"00", X"00", X"0d", X"6e", X"78", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"78", X"56", X"09", X"00", X"00", X"01", X"02", X"03", X"04", X"02", X"00", X"00", X"00", X"01", X"00", X"00", X"02", X"00", X"00", X"01", X"01", X"00", X"02", X"00", X"00", X"00", X"03", X"00", X"00", X"03", X"00", X"00", X"00", X"02", X"00", X"01", X"01", X"00", X"01", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"02", X"00", X"03", X"01", X"02", X"00", X"00", X"09", X"56", X"77", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"79", X"7c", X"7f", X"7e", X"7e", X"77", X"06", X"00", X"00", X"00", X"00", X"00", X"02", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"05", X"01", X"03", X"00", X"00", X"00", X"00", X"03", X"01", X"05", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"01", X"01", X"00", X"00", X"00", X"01", X"00", X"00", X"08", X"74", X"7b", X"7e", X"7f", X"7e", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"78", X"2e", X"00", X"00", X"02", X"00", X"00", X"01", X"02", X"02", X"00", X"00", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"01", X"00", X"00", X"01", X"01", X"00", X"00", X"02", X"00", X"00", X"2d", X"77", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7a", X"68", X"06", X"06", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"02", X"02", X"00", X"02", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"02", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"06", X"67", X"7b", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7c", X"7f", X"7f", X"7f", X"7f", X"7c", X"79", X"7c", X"7c", X"7a", X"74", X"2d", X"04", X"00", X"04", X"02", X"03", X"01", X"00", X"00", X"01", X"02", X"02", X"02", X"01", X"00", X"00", X"00", X"00", X"01", X"02", X"02", X"02", X"01", X"00", X"00", X"00", X"03", X"02", X"02", X"00", X"05", X"2e", X"75", X"7a", X"7e", X"7d", X"7b", X"7c", X"7f", X"7e", X"7d", X"7c", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7b", X"77", X"5b", X"2d", X"12", X"04", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"02", X"02", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"13", X"27", X"53", X"77", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7f", X"7e", X"7f", X"7f", X"7d", X"7d", X"7c", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7d", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7b", X"74", X"3f", X"2c", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"2c", X"3f", X"74", X"7b", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7e", X"7f", X"7b", X"7b", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7e", X"7a", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f"
    );

    constant g_rom : RomType := (
        X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"7f", X"66", X"5b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7f", X"31", X"10", X"0c", X"29", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"1e", X"08", X"0c", X"0b", X"0a", X"11", X"6c", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"73", X"0e", X"0c", X"0b", X"08", X"08", X"0b", X"08", X"0b", X"3b", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"54", X"0c", X"0c", X"08", X"09", X"08", X"08", X"09", X"08", X"0a", X"0b", X"26", X"7f", X"7f", X"7d", X"7c", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"33", X"09", X"0b", X"08", X"0a", X"09", X"08", X"08", X"0b", X"08", X"08", X"0c", X"0a", X"0a", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"29", X"0e", X"0b", X"06", X"09", X"09", X"0b", X"0a", X"09", X"08", X"0a", X"0a", X"08", X"08", X"0b", X"0e", X"66", X"7f", X"7f", X"7e", X"7f", X"7d", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"24", X"0a", X"09", X"09", X"0a", X"08", X"09", X"09", X"09", X"09", X"09", X"0a", X"0a", X"09", X"09", X"08", X"09", X"0e", X"65", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"0d", X"08", X"0b", X"0a", X"09", X"08", X"08", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"0a", X"0a", X"0a", X"09", X"0a", X"55", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7f", X"19", X"0c", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"08", X"08", X"09", X"09", X"08", X"08", X"09", X"0a", X"0a", X"0a", X"08", X"07", X"0c", X"4e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"16", X"0c", X"09", X"09", X"08", X"08", X"08", X"09", X"0a", X"0a", X"09", X"08", X"09", X"09", X"08", X"09", X"09", X"0a", X"0a", X"09", X"0a", X"09", X"09", X"07", X"5d", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"1a", X"09", X"08", X"0a", X"09", X"0a", X"09", X"09", X"08", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"0b", X"0d", X"59", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"2c", X"0e", X"0a", X"09", X"09", X"0a", X"0a", X"0a", X"09", X"09", X"09", X"09", X"09", X"0a", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"0a", X"0a", X"08", X"09", X"0e", X"6e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"32", X"0c", X"08", X"09", X"09", X"09", X"09", X"08", X"09", X"0a", X"0a", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"0a", X"07", X"0a", X"08", X"08", X"0a", X"0a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"57", X"0c", X"0a", X"09", X"0b", X"0a", X"07", X"09", X"09", X"0a", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"08", X"08", X"08", X"09", X"0a", X"09", X"08", X"0b", X"07", X"09", X"0b", X"16", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"73", X"0b", X"09", X"09", X"08", X"07", X"09", X"0a", X"0a", X"08", X"0a", X"0b", X"12", X"29", X"39", X"44", X"4b", X"4c", X"47", X"3b", X"2a", X"15", X"0a", X"0c", X"08", X"09", X"09", X"0b", X"0a", X"09", X"0a", X"08", X"0b", X"21", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"0f", X"09", X"0a", X"09", X"0a", X"07", X"06", X"0c", X"0a", X"0e", X"33", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7e", X"7e", X"7e", X"34", X"0e", X"07", X"0c", X"08", X"07", X"0b", X"08", X"09", X"0a", X"0c", X"44", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"19", X"0b", X"09", X"08", X"09", X"08", X"09", X"0a", X"16", X"70", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"3d", X"6b", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"76", X"15", X"0b", X"0b", X"07", X"08", X"07", X"0a", X"07", X"0b", X"75", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7d", X"7f", X"7f", X"46", X"0c", X"09", X"0a", X"0a", X"08", X"0a", X"12", X"50", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7e", X"7d", X"7f", X"23", X"0a", X"09", X"7f", X"7f", X"7e", X"7c", X"7e", X"7f", X"7f", X"7f", X"51", X"12", X"09", X"0c", X"08", X"08", X"0a", X"0a", X"13", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"0c", X"0b", X"0a", X"08", X"08", X"0c", X"17", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"7f", X"7d", X"7e", X"16", X"0c", X"09", X"0b", X"67", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7d", X"16", X"0b", X"0d", X"0b", X"07", X"0a", X"0a", X"22", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"12", X"0b", X"0b", X"09", X"0b", X"0b", X"2e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"19", X"09", X"0b", X"08", X"0d", X"18", X"7f", X"7f", X"7d", X"7e", X"7d", X"7b", X"7e", X"7e", X"7f", X"7f", X"34", X"09", X"0a", X"09", X"08", X"0b", X"09", X"77", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"46", X"09", X"09", X"07", X"0b", X"0a", X"1c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7d", X"0b", X"0a", X"0b", X"0c", X"0b", X"08", X"0b", X"58", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"1f", X"0e", X"07", X"0b", X"09", X"0c", X"0b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"75", X"0c", X"0a", X"0a", X"07", X"09", X"26", X"7f", X"7e", X"7f", X"7f", X"7f", X"7b", X"7d", X"7f", X"7f", X"6a", X"12", X"08", X"08", X"07", X"08", X"06", X"09", X"0c", X"14", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"2c", X"0c", X"08", X"09", X"09", X"0a", X"41", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"1d", X"0b", X"0b", X"0b", X"0a", X"12", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"5b", X"0f", X"0a", X"07", X"09", X"07", X"08", X"09", X"0c", X"08", X"09", X"6e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"14", X"0c", X"07", X"07", X"0a", X"0d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"4b", X"0b", X"0a", X"09", X"09", X"0c", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"47", X"0f", X"0a", X"0d", X"0c", X"0a", X"09", X"0b", X"0a", X"05", X"09", X"07", X"08", X"7d", X"7e", X"7e", X"7b", X"7c", X"7e", X"7e", X"7f", X"7f", X"7e", X"7f", X"7e", X"0b", X"0a", X"0a", X"0b", X"09", X"17", X"7f", X"7f", X"7e", X"7d", X"7d", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"0a", X"0a", X"05", X"0a", X"0c", X"1b", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"6e", X"6a", X"6d", X"6f", X"2e", X"0d", X"0c", X"15", X"6d", X"71", X"72", X"70", X"70", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"27", X"0b", X"06", X"08", X"08", X"09", X"7b", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7f", X"7f", X"7e", X"7e", X"7f", X"44", X"0b", X"0a", X"0c", X"0c", X"0a", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7e", X"14", X"0c", X"0d", X"52", X"7f", X"7e", X"7e", X"7f", X"7f", X"7e", X"7e", X"7e", X"7c", X"7e", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"08", X"09", X"0b", X"0c", X"0e", X"33", X"7f", X"7c", X"7e", X"7f", X"7d", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7c", X"7d", X"7d", X"7e", X"0c", X"09", X"0a", X"08", X"0d", X"2e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"40", X"0b", X"09", X"09", X"7e", X"7d", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"3d", X"0b", X"09", X"0a", X"09", X"0c", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7c", X"7f", X"7f", X"7f", X"37", X"0a", X"09", X"09", X"0a", X"09", X"71", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"70", X"0c", X"0a", X"0b", X"10", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7c", X"72", X"0b", X"0b", X"0a", X"0a", X"0a", X"2a", X"7f", X"7f", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7e", X"7c", X"7f", X"7f", X"7f", X"7f", X"0e", X"0a", X"08", X"07", X"09", X"08", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"12", X"0b", X"0a", X"0c", X"33", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"5e", X"0c", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"0c", X"0a", X"09", X"0a", X"0b", X"0a", X"7f", X"7e", X"7f", X"7f", X"7d", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"48", X"0b", X"07", X"0a", X"09", X"0a", X"1b", X"7f", X"7e", X"7c", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"25", X"0c", X"0b", X"08", X"0a", X"7b", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"32", X"14", X"09", X"0b", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"22", X"08", X"09", X"07", X"09", X"0c", X"41", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"07", X"09", X"09", X"0a", X"09", X"0a", X"62", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7e", X"7d", X"7f", X"7f", X"7f", X"7e", X"0e", X"08", X"09", X"0a", X"09", X"7e", X"7f", X"7e", X"7e", X"7f", X"54", X"0f", X"0b", X"09", X"0a", X"09", X"08", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"61", X"0a", X"08", X"0a", X"09", X"08", X"0a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"63", X"0a", X"09", X"0a", X"07", X"0b", X"0b", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7d", X"7d", X"7f", X"7f", X"13", X"08", X"0c", X"0c", X"0b", X"23", X"7f", X"7d", X"32", X"13", X"09", X"09", X"09", X"08", X"0a", X"08", X"09", X"09", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"09", X"0c", X"08", X"0a", X"09", X"08", X"69", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"1f", X"09", X"0a", X"0a", X"09", X"0a", X"08", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"56", X"0c", X"09", X"09", X"0b", X"0c", X"12", X"12", X"0b", X"09", X"0a", X"08", X"09", X"0b", X"0a", X"0a", X"09", X"08", X"09", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7e", X"7f", X"7f", X"0c", X"08", X"09", X"09", X"09", X"0a", X"30", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"0b", X"0b", X"08", X"09", X"0b", X"09", X"0b", X"7e", X"7f", X"7e", X"7d", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"18", X"0a", X"09", X"09", X"08", X"06", X"08", X"06", X"0a", X"09", X"09", X"07", X"08", X"08", X"08", X"0a", X"09", X"0a", X"0e", X"7f", X"7f", X"7f", X"7d", X"7e", X"7e", X"7d", X"7f", X"7f", X"7d", X"0f", X"0a", X"09", X"09", X"09", X"0b", X"0b", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7e", X"33", X"0a", X"0a", X"0a", X"0a", X"08", X"09", X"0c", X"7f", X"7e", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"44", X"0b", X"09", X"0a", X"09", X"08", X"0a", X"07", X"0c", X"07", X"09", X"0b", X"25", X"1f", X"0b", X"0c", X"05", X"09", X"0c", X"19", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7e", X"7f", X"0f", X"0a", X"09", X"0a", X"0a", X"0a", X"0a", X"50", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"0f", X"0b", X"0a", X"0d", X"0a", X"09", X"07", X"09", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"07", X"08", X"08", X"09", X"06", X"08", X"0d", X"0c", X"0b", X"0b", X"1b", X"69", X"7f", X"0c", X"0a", X"06", X"0a", X"0b", X"0b", X"2a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7e", X"0d", X"07", X"0b", X"09", X"0a", X"09", X"0c", X"15", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"09", X"0a", X"06", X"08", X"08", X"0b", X"0a", X"0b", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"4d", X"0b", X"09", X"0a", X"06", X"0a", X"0a", X"09", X"0c", X"0e", X"4f", X"7f", X"7c", X"7f", X"0c", X"08", X"0b", X"09", X"09", X"0a", X"44", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"0b", X"0b", X"09", X"08", X"09", X"0a", X"0a", X"0e", X"7d", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"53", X"0b", X"08", X"0b", X"0a", X"0a", X"08", X"08", X"07", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"0f", X"07", X"09", X"0a", X"0a", X"09", X"0a", X"10", X"5d", X"7f", X"7e", X"7f", X"7f", X"55", X"0a", X"0b", X"09", X"09", X"0a", X"0c", X"5d", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"08", X"09", X"09", X"0a", X"0a", X"0a", X"08", X"0b", X"7b", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"15", X"07", X"09", X"07", X"0b", X"09", X"0b", X"08", X"08", X"4f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"4f", X"0a", X"0a", X"09", X"08", X"0e", X"27", X"63", X"7f", X"7f", X"7c", X"7e", X"7f", X"7f", X"24", X"0a", X"08", X"08", X"08", X"09", X"0a", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"53", X"0c", X"09", X"07", X"09", X"09", X"09", X"08", X"08", X"42", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"09", X"0a", X"09", X"0b", X"08", X"09", X"08", X"09", X"0b", X"15", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"1a", X"0c", X"0b", X"09", X"48", X"7f", X"7d", X"7f", X"7e", X"7f", X"7f", X"7e", X"7f", X"7d", X"0c", X"0b", X"09", X"08", X"0b", X"09", X"0a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7d", X"7f", X"7f", X"16", X"0a", X"09", X"09", X"09", X"08", X"08", X"08", X"0b", X"0b", X"7f", X"7e", X"7f", X"7f", X"7f", X"6b", X"0a", X"0c", X"0a", X"0a", X"09", X"09", X"0a", X"0a", X"08", X"0b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"3d", X"65", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"1e", X"0b", X"05", X"09", X"0b", X"07", X"0b", X"11", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7d", X"7f", X"0e", X"09", X"08", X"0a", X"09", X"09", X"0b", X"09", X"08", X"0b", X"7f", X"7f", X"7d", X"7f", X"7f", X"43", X"0d", X"09", X"09", X"09", X"0a", X"0a", X"09", X"07", X"0b", X"09", X"66", X"7f", X"7e", X"7f", X"7e", X"7d", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7e", X"09", X"07", X"0b", X"09", X"08", X"0a", X"0c", X"1f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"6e", X"0a", X"09", X"09", X"09", X"0a", X"0a", X"09", X"07", X"0d", X"0d", X"6d", X"7d", X"7d", X"7e", X"7f", X"27", X"0b", X"0a", X"09", X"0b", X"09", X"0a", X"09", X"07", X"09", X"0b", X"24", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"1f", X"0c", X"0b", X"08", X"08", X"05", X"0b", X"08", X"2e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"2b", X"0d", X"0a", X"0a", X"09", X"08", X"07", X"0c", X"09", X"0b", X"0c", X"44", X"7e", X"7c", X"7f", X"7f", X"19", X"0c", X"0b", X"09", X"08", X"09", X"09", X"0a", X"09", X"07", X"09", X"0d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7c", X"7f", X"7e", X"7e", X"7f", X"62", X"09", X"09", X"08", X"09", X"0a", X"0b", X"0b", X"0c", X"58", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"0b", X"09", X"07", X"08", X"0c", X"09", X"08", X"0a", X"0a", X"09", X"0e", X"30", X"7b", X"7d", X"7f", X"7f", X"0c", X"0a", X"08", X"09", X"06", X"0a", X"0b", X"08", X"08", X"0a", X"07", X"08", X"17", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"13", X"0b", X"0a", X"0b", X"06", X"09", X"0a", X"09", X"09", X"7c", X"7f", X"7e", X"7f", X"7d", X"7e", X"7e", X"7e", X"7f", X"17", X"0a", X"0b", X"0a", X"09", X"09", X"09", X"0a", X"07", X"09", X"0b", X"0b", X"1a", X"7f", X"7f", X"7f", X"7f", X"09", X"0a", X"08", X"09", X"09", X"08", X"0a", X"0c", X"08", X"0a", X"08", X"0a", X"0c", X"59", X"7f", X"7f", X"7e", X"7f", X"7f", X"7d", X"7e", X"7d", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"2b", X"0e", X"09", X"09", X"07", X"0a", X"09", X"0a", X"0c", X"15", X"7f", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"6b", X"0a", X"09", X"08", X"08", X"0b", X"08", X"09", X"09", X"08", X"0a", X"0b", X"09", X"0f", X"7f", X"7f", X"7f", X"77", X"09", X"09", X"0a", X"09", X"0b", X"09", X"08", X"08", X"09", X"09", X"09", X"09", X"08", X"09", X"7c", X"7f", X"7e", X"7f", X"7f", X"7f", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"68", X"08", X"0a", X"0a", X"09", X"07", X"0b", X"06", X"0b", X"0b", X"3f", X"7f", X"7f", X"7e", X"7e", X"7d", X"7d", X"7f", X"7f", X"09", X"09", X"09", X"0a", X"0a", X"09", X"08", X"08", X"0a", X"08", X"0a", X"0a", X"09", X"09", X"7d", X"7e", X"7f", X"49", X"0a", X"0a", X"09", X"0a", X"07", X"09", X"08", X"09", X"0a", X"0a", X"0a", X"09", X"09", X"0a", X"1a", X"7f", X"7f", X"7f", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"0b", X"09", X"09", X"08", X"07", X"0b", X"08", X"09", X"0a", X"09", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"18", X"0a", X"09", X"09", X"09", X"0a", X"0a", X"08", X"08", X"07", X"0d", X"0a", X"09", X"07", X"08", X"7c", X"7f", X"7f", X"35", X"0a", X"07", X"09", X"0a", X"09", X"09", X"0a", X"0a", X"09", X"09", X"09", X"09", X"09", X"0a", X"09", X"17", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7d", X"16", X"0c", X"08", X"07", X"0a", X"0a", X"07", X"0a", X"0d", X"0a", X"0b", X"7e", X"7f", X"7e", X"7d", X"7f", X"7d", X"7f", X"1d", X"0e", X"0b", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"0a", X"09", X"0c", X"08", X"62", X"7f", X"7f", X"22", X"0b", X"09", X"09", X"06", X"08", X"0a", X"0a", X"0a", X"09", X"08", X"08", X"08", X"09", X"08", X"08", X"07", X"17", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7e", X"7f", X"1c", X"0a", X"09", X"0a", X"0a", X"07", X"0a", X"09", X"09", X"06", X"09", X"34", X"7f", X"7e", X"7e", X"7e", X"7d", X"7f", X"17", X"08", X"0a", X"09", X"0a", X"0a", X"0a", X"08", X"08", X"09", X"0a", X"09", X"0a", X"08", X"07", X"0a", X"0d", X"45", X"7f", X"7f", X"14", X"0b", X"08", X"09", X"0a", X"08", X"08", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"09", X"0a", X"0a", X"09", X"11", X"71", X"7f", X"7d", X"7e", X"7d", X"7f", X"23", X"0e", X"0c", X"09", X"07", X"09", X"0a", X"0a", X"09", X"0b", X"0a", X"0c", X"7e", X"7e", X"7f", X"7f", X"7f", X"71", X"12", X"09", X"07", X"09", X"09", X"0a", X"09", X"09", X"09", X"09", X"09", X"09", X"07", X"0b", X"08", X"08", X"09", X"09", X"27", X"7f", X"7f", X"0b", X"0c", X"08", X"0a", X"09", X"09", X"0a", X"08", X"08", X"09", X"0a", X"0a", X"09", X"09", X"09", X"07", X"08", X"0b", X"0c", X"0c", X"3c", X"7f", X"7f", X"7f", X"12", X"0b", X"07", X"09", X"0a", X"08", X"09", X"07", X"08", X"08", X"0b", X"0b", X"35", X"7f", X"7e", X"7f", X"7f", X"3b", X"0b", X"07", X"09", X"0b", X"0b", X"09", X"09", X"09", X"09", X"0a", X"0a", X"09", X"08", X"09", X"07", X"09", X"0c", X"08", X"0b", X"14", X"7f", X"7f", X"7f", X"19", X"08", X"0b", X"0c", X"09", X"09", X"08", X"08", X"09", X"0a", X"0a", X"0a", X"09", X"09", X"09", X"09", X"0a", X"0b", X"0c", X"0a", X"0b", X"35", X"7f", X"4d", X"09", X"0a", X"08", X"08", X"0b", X"09", X"09", X"0c", X"09", X"08", X"0a", X"7c", X"7f", X"7f", X"37", X"0b", X"08", X"0c", X"0a", X"0b", X"0a", X"08", X"08", X"09", X"0a", X"0b", X"09", X"09", X"08", X"08", X"08", X"0b", X"09", X"0a", X"0c", X"18", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"1d", X"0a", X"09", X"08", X"08", X"08", X"09", X"09", X"09", X"09", X"08", X"08", X"09", X"0a", X"09", X"07", X"08", X"08", X"07", X"09", X"0f", X"2c", X"42", X"38", X"34", X"13", X"08", X"0a", X"0b", X"07", X"09", X"0b", X"16", X"51", X"2a", X"0d", X"0b", X"0b", X"0a", X"09", X"0a", X"0a", X"07", X"09", X"08", X"08", X"09", X"09", X"09", X"0a", X"0a", X"09", X"09", X"08", X"0b", X"1d", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"67", X"1f", X"0d", X"0b", X"09", X"08", X"07", X"08", X"08", X"09", X"09", X"09", X"0a", X"09", X"0a", X"0b", X"08", X"07", X"09", X"0a", X"09", X"09", X"07", X"0d", X"0f", X"21", X"22", X"22", X"21", X"0f", X"0d", X"07", X"09", X"09", X"0a", X"09", X"06", X"0a", X"0b", X"09", X"09", X"09", X"09", X"0a", X"0a", X"0a", X"06", X"07", X"07", X"09", X"0b", X"0c", X"1e", X"67", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7e", X"7e", X"7e", X"17", X"0d", X"09", X"09", X"0a", X"09", X"0b", X"07", X"08", X"06", X"09", X"0a", X"08", X"09", X"0a", X"0b", X"0a", X"0c", X"09", X"0b", X"05", X"08", X"09", X"09", X"09", X"09", X"07", X"05", X"0a", X"08", X"0b", X"0a", X"0a", X"0a", X"08", X"08", X"0a", X"0a", X"08", X"09", X"08", X"09", X"06", X"0b", X"0a", X"0b", X"0d", X"1f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7d", X"7e", X"7f", X"42", X"15", X"09", X"0b", X"09", X"0b", X"09", X"09", X"0c", X"0a", X"0a", X"0b", X"08", X"07", X"09", X"08", X"0b", X"0a", X"0b", X"09", X"0a", X"08", X"08", X"0a", X"09", X"0b", X"0a", X"0b", X"08", X"09", X"0a", X"08", X"09", X"0a", X"0a", X"08", X"08", X"09", X"0a", X"0a", X"0b", X"09", X"13", X"42", X"7d", X"7f", X"7d", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7c", X"7f", X"7c", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7a", X"19", X"10", X"09", X"0a", X"07", X"0b", X"0a", X"08", X"09", X"09", X"0c", X"09", X"07", X"09", X"07", X"08", X"0a", X"09", X"0a", X"0a", X"09", X"0a", X"08", X"07", X"0a", X"07", X"0a", X"09", X"0a", X"0b", X"0a", X"0b", X"0c", X"09", X"09", X"09", X"10", X"1b", X"79", X"7f", X"7e", X"7d", X"7e", X"7e", X"7d", X"7f", X"7f", X"7b", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"3d", X"15", X"07", X"0b", X"09", X"0a", X"0a", X"08", X"09", X"0a", X"09", X"08", X"08", X"09", X"0a", X"09", X"09", X"0a", X"09", X"09", X"08", X"09", X"0b", X"09", X"09", X"09", X"09", X"08", X"0a", X"06", X"15", X"3e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"6c", X"44", X"2c", X"1c", X"0e", X"0a", X"0b", X"0a", X"09", X"0a", X"0a", X"0a", X"0a", X"09", X"09", X"09", X"0a", X"08", X"09", X"0a", X"0a", X"0e", X"1d", X"2c", X"3e", X"64", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7c", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7c", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7d", X"7c", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"55", X"49", X"2d", X"18", X"16", X"0b", X"0a", X"16", X"17", X"2d", X"48", X"55", X"7e", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7c", X"7d", X"7c", X"7f", X"7f", X"7e", X"7f", X"7e", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"7d", X"7e", X"7e", X"7d", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f"
    );

    constant b_rom : RomType := (
        X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7e", X"7e", X"7d", X"7d", X"7f", X"7f", X"7f", X"7c", X"7c", X"7d", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"72", X"68", X"7f", X"7f", X"7d", X"7d", X"7d", X"7e", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7e", X"7e", X"7d", X"7c", X"7f", X"7f", X"7f", X"7f", X"44", X"2a", X"2b", X"41", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7d", X"7d", X"7d", X"7e", X"7e", X"7d", X"7f", X"7f", X"34", X"25", X"2d", X"2e", X"2a", X"2c", X"7d", X"7f", X"7d", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"27", X"2d", X"2f", X"2c", X"29", X"2d", X"2e", X"2c", X"4d", X"7f", X"7f", X"7d", X"7d", X"7c", X"7e", X"7c", X"7b", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"67", X"27", X"2c", X"2a", X"2d", X"2c", X"2b", X"2b", X"2b", X"2d", X"2e", X"40", X"7f", X"7e", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"47", X"28", X"2f", X"2b", X"2b", X"2b", X"2b", X"2b", X"2e", X"2b", X"2c", X"30", X"2a", X"23", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7b", X"7d", X"7f", X"3e", X"2d", X"2f", X"2c", X"2d", X"2a", X"2b", X"2a", X"2c", X"2c", X"2e", X"2d", X"2a", X"29", X"2d", X"29", X"72", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7a", X"7e", X"7f", X"7f", X"38", X"2b", X"2f", X"2a", X"29", X"2d", X"2d", X"2b", X"2a", X"2a", X"2a", X"2a", X"2a", X"2c", X"2c", X"2d", X"2b", X"29", X"77", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"27", X"2a", X"2b", X"2a", X"2a", X"2b", X"2e", X"2e", X"2d", X"2c", X"2b", X"2b", X"2d", X"2d", X"2c", X"2c", X"2c", X"2b", X"29", X"25", X"67", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"2d", X"2d", X"2f", X"2c", X"2b", X"2d", X"2c", X"2c", X"2c", X"2e", X"2e", X"2d", X"2d", X"2e", X"2e", X"2c", X"2b", X"2c", X"2c", X"2b", X"29", X"29", X"61", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"33", X"31", X"2a", X"2a", X"2c", X"2d", X"2f", X"2d", X"29", X"29", X"2d", X"2e", X"2e", X"2d", X"2e", X"2d", X"2b", X"2a", X"2b", X"2c", X"2f", X"2f", X"2d", X"24", X"6c", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7a", X"7f", X"7f", X"2e", X"2a", X"2c", X"2e", X"2c", X"2b", X"2c", X"2d", X"2d", X"2b", X"2a", X"2b", X"2c", X"2d", X"2d", X"2b", X"2a", X"2a", X"2a", X"2b", X"2c", X"2e", X"2e", X"2d", X"2b", X"27", X"69", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"45", X"2e", X"2c", X"2a", X"2c", X"2c", X"2b", X"2a", X"2c", X"2c", X"2d", X"2c", X"2a", X"2a", X"2d", X"2c", X"2a", X"28", X"2a", X"2a", X"2c", X"2d", X"2d", X"2e", X"2b", X"29", X"2b", X"2a", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"46", X"2a", X"2b", X"2e", X"2b", X"2a", X"29", X"2c", X"2d", X"2d", X"2d", X"2d", X"2d", X"2c", X"2c", X"2d", X"2c", X"2a", X"2a", X"2b", X"2c", X"2e", X"2d", X"2d", X"29", X"2c", X"2b", X"2c", X"2b", X"23", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"6d", X"2a", X"2b", X"2b", X"2d", X"2d", X"2b", X"2c", X"2d", X"2d", X"2d", X"2d", X"2e", X"2e", X"2e", X"2e", X"2d", X"2d", X"2c", X"2c", X"2e", X"2e", X"2f", X"2d", X"2c", X"2b", X"2d", X"31", X"29", X"29", X"2b", X"2d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7b", X"7e", X"7f", X"7f", X"7d", X"23", X"28", X"2d", X"2d", X"2e", X"2e", X"2e", X"2b", X"2a", X"2c", X"30", X"35", X"45", X"51", X"5c", X"62", X"62", X"5e", X"58", X"49", X"35", X"2c", X"2d", X"2a", X"2f", X"2c", X"2a", X"28", X"2a", X"2c", X"2a", X"28", X"38", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"25", X"29", X"30", X"2d", X"2f", X"2c", X"2b", X"32", X"2d", X"2e", X"48", X"7f", X"7d", X"7d", X"7e", X"7d", X"7c", X"79", X"79", X"7d", X"7e", X"7f", X"7f", X"49", X"2b", X"29", X"30", X"2c", X"2b", X"30", X"2d", X"2d", X"2b", X"28", X"57", X"7f", X"7d", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7e", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"31", X"2b", X"28", X"28", X"2d", X"2c", X"2d", X"2a", X"2d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"50", X"7e", X"7f", X"7d", X"7f", X"7f", X"7c", X"7f", X"7f", X"2f", X"28", X"2c", X"2c", X"2e", X"2c", X"2e", X"2a", X"26", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7e", X"7e", X"7d", X"7d", X"7e", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"55", X"2a", X"2f", X"30", X"2e", X"2a", X"28", X"31", X"65", X"7f", X"7c", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"39", X"27", X"22", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"65", X"2e", X"29", X"2e", X"2d", X"2e", X"31", X"29", X"27", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"24", X"2b", X"2d", X"2a", X"2a", X"31", X"32", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7c", X"7f", X"2c", X"2c", X"2d", X"28", X"72", X"7f", X"7f", X"7f", X"7f", X"7d", X"7b", X"79", X"7d", X"7f", X"2f", X"29", X"2a", X"29", X"2b", X"2d", X"28", X"35", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"29", X"2a", X"2c", X"2a", X"2e", X"2a", X"47", X"7f", X"7f", X"7a", X"79", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"2d", X"25", X"2a", X"2a", X"2a", X"2a", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"49", X"29", X"2d", X"2c", X"2a", X"31", X"27", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7d", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"56", X"26", X"2b", X"2a", X"2e", X"2e", X"37", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"27", X"2d", X"2b", X"2b", X"2a", X"25", X"26", X"6b", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7b", X"7c", X"7f", X"38", X"2f", X"29", X"2d", X"2e", X"2c", X"21", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"23", X"29", X"2d", X"2c", X"29", X"39", X"7f", X"7f", X"7d", X"7d", X"7d", X"7f", X"7f", X"7d", X"7f", X"76", X"29", X"27", X"2c", X"2e", X"31", X"33", X"32", X"2f", X"29", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"3f", X"29", X"2a", X"2a", X"29", X"27", X"56", X"7f", X"7d", X"7d", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7e", X"7c", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"37", X"2a", X"2a", X"29", X"2b", X"2d", X"7f", X"7f", X"7e", X"7d", X"7e", X"7e", X"7f", X"7f", X"7f", X"6a", X"28", X"2b", X"2e", X"31", X"2a", X"28", X"29", X"2b", X"2b", X"25", X"7d", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"2c", X"2b", X"29", X"2b", X"30", X"2a", X"7f", X"7f", X"7f", X"7d", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7d", X"7d", X"7d", X"7d", X"7f", X"7f", X"5d", X"2b", X"2f", X"2c", X"27", X"24", X"7f", X"7f", X"7d", X"7d", X"7d", X"7f", X"7e", X"7c", X"7f", X"5e", X"31", X"29", X"2b", X"2c", X"2b", X"2c", X"2e", X"30", X"2b", X"31", X"2b", X"22", X"7f", X"7f", X"7d", X"7f", X"7f", X"7e", X"7c", X"7d", X"7c", X"7d", X"7f", X"7f", X"20", X"28", X"2e", X"32", X"2c", X"2c", X"7f", X"7f", X"7b", X"7c", X"7e", X"7f", X"7e", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"1d", X"25", X"26", X"2c", X"2a", X"31", X"7f", X"7f", X"7e", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"49", X"2d", X"2f", X"33", X"7f", X"7f", X"7f", X"7a", X"77", X"7f", X"7f", X"7e", X"7d", X"7b", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"37", X"29", X"2a", X"2c", X"27", X"1d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7b", X"7d", X"7d", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"5d", X"2b", X"2a", X"2d", X"2e", X"25", X"7f", X"7e", X"7f", X"7f", X"7f", X"7e", X"7c", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"2f", X"2c", X"28", X"65", X"7f", X"7f", X"7d", X"7c", X"7e", X"7d", X"7d", X"7d", X"7f", X"7f", X"7f", X"7d", X"7f", X"7d", X"7f", X"7f", X"7d", X"7f", X"24", X"2d", X"2c", X"2c", X"2d", X"4a", X"7f", X"7e", X"7f", X"7f", X"7f", X"7c", X"7c", X"7b", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"26", X"2a", X"2b", X"29", X"2d", X"46", X"7f", X"7e", X"7f", X"7f", X"7e", X"7d", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"4c", X"27", X"27", X"1e", X"7f", X"7f", X"7f", X"7c", X"7c", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7b", X"7e", X"7f", X"55", X"2b", X"28", X"2a", X"29", X"24", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"79", X"7b", X"7f", X"7f", X"7f", X"7f", X"7f", X"4a", X"28", X"2c", X"2c", X"2a", X"24", X"7f", X"7f", X"7d", X"7e", X"7f", X"7e", X"7e", X"7f", X"7f", X"7d", X"7d", X"7d", X"7f", X"7f", X"27", X"2a", X"29", X"28", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7b", X"7d", X"7f", X"7f", X"7d", X"7c", X"7f", X"7f", X"7f", X"24", X"28", X"29", X"2b", X"26", X"3e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7c", X"7f", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"23", X"2b", X"2e", X"2e", X"2b", X"24", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"2b", X"2d", X"2d", X"2a", X"49", X"7f", X"7f", X"7c", X"7f", X"7f", X"7f", X"7f", X"7c", X"7f", X"77", X"23", X"7f", X"78", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"23", X"28", X"2b", X"2f", X"2c", X"22", X"7f", X"7f", X"7d", X"7e", X"7e", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7e", X"7f", X"5a", X"28", X"28", X"2d", X"2e", X"2a", X"2e", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"3c", X"28", X"2b", X"2b", X"24", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"4b", X"36", X"2f", X"27", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"31", X"26", X"2e", X"2d", X"2d", X"2d", X"59", X"7f", X"7e", X"7f", X"7f", X"7b", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"23", X"2d", X"2c", X"2b", X"29", X"23", X"6f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"20", X"25", X"2d", X"2f", X"24", X"7f", X"7d", X"7f", X"7f", X"7f", X"64", X"2d", X"30", X"2e", X"2e", X"2d", X"23", X"7f", X"7e", X"7f", X"7f", X"7e", X"7d", X"7e", X"7f", X"7f", X"6d", X"22", X"28", X"2c", X"2d", X"2c", X"26", X"7f", X"7f", X"7f", X"7f", X"7e", X"7c", X"7f", X"7f", X"7d", X"7f", X"7f", X"72", X"26", X"2b", X"2d", X"2a", X"30", X"27", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7f", X"7f", X"7f", X"7f", X"2f", X"2f", X"33", X"30", X"2b", X"3a", X"7f", X"7f", X"47", X"30", X"29", X"28", X"25", X"25", X"2c", X"2c", X"30", X"26", X"7f", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"21", X"2b", X"2b", X"2e", X"2d", X"25", X"76", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7d", X"7f", X"7f", X"33", X"28", X"2d", X"2d", X"2c", X"2e", X"24", X"7f", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"66", X"28", X"2c", X"2c", X"2d", X"2f", X"33", X"33", X"2c", X"2c", X"30", X"2f", X"2c", X"27", X"26", X"2d", X"30", X"2e", X"24", X"7f", X"7c", X"7c", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"25", X"28", X"2b", X"2c", X"2c", X"27", X"42", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"24", X"2c", X"2c", X"2d", X"2d", X"2c", X"25", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7d", X"7c", X"7d", X"7f", X"7f", X"27", X"23", X"27", X"2a", X"2c", X"2f", X"31", X"2c", X"2d", X"29", X"29", X"2e", X"2f", X"2c", X"2c", X"30", X"2d", X"2c", X"24", X"7f", X"7b", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"29", X"2d", X"2b", X"2a", X"2b", X"29", X"22", X"7f", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"47", X"25", X"2c", X"2e", X"2e", X"2c", X"2d", X"27", X"7f", X"7e", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"5a", X"29", X"29", X"2b", X"2d", X"2b", X"2b", X"27", X"2b", X"29", X"2f", X"30", X"43", X"3d", X"2f", X"33", X"2a", X"2c", X"2d", X"30", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"2a", X"2d", X"2c", X"2c", X"2c", X"29", X"26", X"64", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"28", X"2c", X"2c", X"2f", X"2c", X"2c", X"2c", X"24", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"25", X"2f", X"2f", X"31", X"31", X"30", X"2e", X"29", X"2d", X"2a", X"34", X"7d", X"7f", X"23", X"2b", X"2a", X"2d", X"2d", X"2f", X"44", X"7f", X"7e", X"7f", X"7f", X"7d", X"7d", X"7e", X"7d", X"7e", X"7f", X"27", X"2a", X"2d", X"2c", X"2c", X"2b", X"2b", X"2c", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"25", X"2e", X"29", X"2a", X"2a", X"2e", X"2b", X"24", X"7f", X"7f", X"7f", X"7e", X"7e", X"7d", X"7d", X"7f", X"7f", X"5d", X"28", X"2d", X"30", X"2b", X"2a", X"2a", X"2c", X"2f", X"2f", X"68", X"7f", X"7f", X"7f", X"20", X"24", X"2d", X"2c", X"2c", X"2b", X"5c", X"7f", X"7c", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"25", X"2e", X"2d", X"2c", X"2c", X"2c", X"2d", X"27", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"60", X"25", X"2a", X"2d", X"2d", X"2d", X"2a", X"2a", X"20", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"26", X"27", X"2c", X"2b", X"2a", X"2a", X"2b", X"30", X"75", X"7f", X"7d", X"7f", X"7f", X"6c", X"2a", X"2d", X"2b", X"2b", X"29", X"27", X"6f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"22", X"2b", X"2d", X"2d", X"2d", X"2d", X"2d", X"26", X"7f", X"7e", X"7d", X"7e", X"7d", X"7f", X"7f", X"2b", X"28", X"2d", X"2a", X"2d", X"2c", X"2d", X"2a", X"23", X"5f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"67", X"2b", X"2c", X"2e", X"2c", X"30", X"45", X"77", X"7f", X"7b", X"7c", X"7e", X"7c", X"7f", X"3e", X"2e", X"2d", X"2d", X"2c", X"27", X"1b", X"7f", X"7f", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"5e", X"29", X"2d", X"2a", X"2b", X"2a", X"2c", X"2f", X"29", X"55", X"7f", X"7f", X"7f", X"7c", X"7f", X"7f", X"22", X"29", X"2a", X"2d", X"2a", X"2e", X"2c", X"2b", X"26", X"29", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7f", X"31", X"2d", X"2d", X"24", X"59", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7f", X"28", X"30", X"2e", X"2a", X"2d", X"25", X"1e", X"7f", X"7f", X"7e", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"26", X"27", X"2b", X"2d", X"2d", X"2b", X"2b", X"2c", X"29", X"1d", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"26", X"2a", X"2a", X"2c", X"2c", X"2e", X"2e", X"2d", X"28", X"25", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"4e", X"75", X"7f", X"7f", X"7f", X"7f", X"7e", X"7c", X"7d", X"7d", X"7e", X"7f", X"7f", X"2d", X"29", X"2a", X"2d", X"2f", X"2a", X"28", X"28", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"23", X"26", X"2b", X"2d", X"2d", X"2e", X"2d", X"2a", X"22", X"1e", X"7f", X"7f", X"7f", X"7e", X"7f", X"5a", X"2d", X"29", X"2a", X"29", X"2c", X"2e", X"2e", X"2d", X"2d", X"26", X"78", X"7f", X"7b", X"7f", X"7f", X"7f", X"7f", X"7d", X"7b", X"79", X"7c", X"7f", X"7f", X"7f", X"7e", X"7b", X"7c", X"7e", X"7f", X"7f", X"25", X"28", X"2f", X"2c", X"2a", X"2a", X"27", X"35", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7d", X"7b", X"7f", X"7f", X"25", X"29", X"2b", X"2e", X"2f", X"2e", X"2c", X"28", X"2a", X"24", X"7d", X"7f", X"7f", X"7d", X"7f", X"3f", X"2c", X"2b", X"2a", X"2b", X"2a", X"2f", X"2f", X"2e", X"2d", X"2c", X"3a", X"7f", X"7d", X"7c", X"7d", X"7f", X"7f", X"7d", X"7c", X"7f", X"7e", X"7a", X"7a", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"34", X"29", X"2b", X"2a", X"2c", X"29", X"2f", X"26", X"42", X"7f", X"7f", X"7e", X"7e", X"7e", X"7f", X"7e", X"7d", X"7f", X"41", X"2c", X"2d", X"2e", X"2b", X"2a", X"2a", X"2e", X"2b", X"2c", X"2a", X"5b", X"7f", X"7f", X"7e", X"7f", X"31", X"2c", X"2e", X"2c", X"2b", X"2b", X"2a", X"2d", X"2e", X"2c", X"2e", X"29", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7a", X"7b", X"7f", X"74", X"28", X"2e", X"2b", X"2b", X"2d", X"2d", X"2c", X"26", X"66", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"25", X"2a", X"2b", X"2c", X"2f", X"2b", X"2a", X"2c", X"2e", X"2d", X"30", X"4a", X"7f", X"7f", X"7e", X"7f", X"26", X"2d", X"2c", X"2b", X"29", X"2b", X"2d", X"2a", X"2c", X"2e", X"2d", X"27", X"2c", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7c", X"7e", X"7e", X"7f", X"7f", X"7f", X"27", X"29", X"2c", X"2e", X"29", X"2c", X"2c", X"2a", X"23", X"7f", X"7f", X"7f", X"7f", X"7d", X"7e", X"7f", X"7f", X"7f", X"2d", X"27", X"2c", X"2d", X"2d", X"2e", X"2d", X"2c", X"29", X"2a", X"2e", X"2f", X"34", X"7f", X"7f", X"7e", X"7f", X"22", X"2c", X"2d", X"2f", X"2c", X"2a", X"2a", X"2c", X"2a", X"2e", X"2f", X"2d", X"24", X"68", X"7f", X"7e", X"7b", X"7d", X"7d", X"7d", X"7f", X"7d", X"7d", X"7d", X"7c", X"7e", X"7d", X"7f", X"45", X"31", X"2d", X"2c", X"2b", X"2d", X"2b", X"2c", X"2c", X"2c", X"7f", X"7d", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"27", X"29", X"2a", X"2a", X"2e", X"2f", X"2f", X"2c", X"29", X"2a", X"2c", X"2c", X"2a", X"7f", X"7d", X"7f", X"7f", X"28", X"30", X"2d", X"2b", X"2d", X"2c", X"2f", X"2f", X"2a", X"2a", X"2d", X"2f", X"2e", X"25", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"79", X"25", X"2c", X"2e", X"2d", X"2b", X"2f", X"2a", X"2d", X"2b", X"53", X"7f", X"7b", X"7c", X"7f", X"7f", X"7f", X"7f", X"7f", X"22", X"2b", X"2e", X"2d", X"29", X"29", X"2e", X"2f", X"2f", X"2b", X"2d", X"2e", X"2f", X"26", X"7f", X"7d", X"7f", X"5a", X"27", X"2c", X"2b", X"2d", X"2c", X"2e", X"2e", X"2c", X"28", X"27", X"29", X"2b", X"2c", X"28", X"2d", X"7f", X"7f", X"7e", X"7c", X"7f", X"7d", X"7d", X"7f", X"7f", X"7e", X"7f", X"7f", X"21", X"2a", X"2e", X"2d", X"2b", X"2d", X"29", X"27", X"26", X"23", X"7f", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"2d", X"28", X"2c", X"2c", X"2c", X"2b", X"2c", X"2d", X"2d", X"28", X"2e", X"2c", X"2c", X"2b", X"23", X"7f", X"7f", X"7f", X"49", X"2a", X"2d", X"2d", X"2c", X"2a", X"2a", X"2b", X"2b", X"2a", X"2a", X"2c", X"2c", X"2b", X"2b", X"2b", X"2f", X"7f", X"7a", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"2f", X"2e", X"2a", X"29", X"2c", X"2d", X"27", X"29", X"2f", X"28", X"1f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7f", X"36", X"2d", X"2b", X"2b", X"2f", X"2f", X"2c", X"2a", X"2a", X"2a", X"2b", X"2b", X"2c", X"2b", X"2d", X"22", X"71", X"7f", X"7f", X"35", X"29", X"2c", X"2f", X"2a", X"2a", X"29", X"29", X"2b", X"2e", X"2f", X"31", X"2f", X"2d", X"2c", X"2f", X"29", X"2b", X"7f", X"7f", X"7d", X"7c", X"7e", X"7f", X"7f", X"7f", X"2b", X"27", X"2d", X"2f", X"2d", X"2a", X"2d", X"2f", X"2d", X"27", X"24", X"43", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"2c", X"24", X"2a", X"2a", X"2b", X"2d", X"2d", X"2d", X"2c", X"2c", X"2a", X"2a", X"2b", X"2c", X"2b", X"2d", X"29", X"58", X"7f", X"7f", X"2c", X"25", X"26", X"2d", X"30", X"2d", X"2c", X"2c", X"2c", X"2d", X"2e", X"2e", X"2d", X"2d", X"2c", X"2d", X"2e", X"2e", X"2e", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"3b", X"2c", X"2d", X"2c", X"2b", X"2d", X"2d", X"2d", X"2c", X"2f", X"2f", X"28", X"7f", X"7f", X"7f", X"7f", X"7f", X"7a", X"2d", X"2c", X"2a", X"2a", X"2a", X"2a", X"2c", X"2c", X"2e", X"2d", X"2b", X"2b", X"2b", X"30", X"2f", X"2e", X"2b", X"26", X"3d", X"7f", X"7f", X"20", X"2e", X"2f", X"2d", X"2b", X"2b", X"2e", X"2f", X"2f", X"2a", X"29", X"2a", X"2a", X"29", X"29", X"2a", X"2a", X"2e", X"2c", X"2a", X"4f", X"7f", X"7f", X"7f", X"28", X"2c", X"2d", X"2e", X"2e", X"2c", X"2d", X"2e", X"2c", X"29", X"27", X"27", X"4b", X"7f", X"7f", X"7c", X"7f", X"50", X"2b", X"2d", X"31", X"30", X"2e", X"2c", X"2b", X"2d", X"2c", X"29", X"29", X"2d", X"2f", X"30", X"2d", X"2c", X"2e", X"2a", X"27", X"26", X"7f", X"7e", X"7f", X"33", X"2a", X"2b", X"2c", X"29", X"2b", X"2e", X"2e", X"2b", X"2b", X"2d", X"2c", X"2a", X"2a", X"2d", X"2d", X"2a", X"28", X"2b", X"29", X"2c", X"50", X"7f", X"5e", X"2a", X"31", X"2f", X"2d", X"2c", X"29", X"2c", X"31", X"2f", X"2a", X"23", X"7f", X"7f", X"7f", X"4f", X"2f", X"30", X"32", X"2c", X"2b", X"2d", X"2c", X"2f", X"2e", X"2b", X"28", X"28", X"2a", X"31", X"32", X"2d", X"2d", X"27", X"28", X"2b", X"30", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"38", X"30", X"32", X"2d", X"28", X"27", X"2f", X"30", X"2f", X"2f", X"2f", X"2e", X"2c", X"2c", X"2d", X"2a", X"2b", X"2d", X"31", X"31", X"2e", X"45", X"58", X"4f", X"52", X"35", X"29", X"2b", X"2b", X"27", X"28", X"29", X"34", X"6e", X"4b", X"2f", X"2b", X"2b", X"29", X"28", X"27", X"29", X"2b", X"2f", X"2e", X"2e", X"2d", X"2d", X"2e", X"2b", X"26", X"27", X"30", X"32", X"33", X"39", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"75", X"38", X"2c", X"2b", X"2c", X"2d", X"2e", X"30", X"2e", X"2d", X"2b", X"2b", X"2b", X"2b", X"2c", X"30", X"2f", X"2f", X"31", X"2f", X"2b", X"29", X"26", X"2c", X"2e", X"40", X"42", X"41", X"40", X"2e", X"2b", X"26", X"28", X"2c", X"2f", X"31", X"2e", X"30", X"2f", X"2a", X"2a", X"2a", X"2a", X"2c", X"2d", X"31", X"2d", X"2f", X"2b", X"2b", X"28", X"2a", X"36", X"75", X"7f", X"7f", X"7f", X"7f", X"7f", X"7b", X"7c", X"7c", X"7f", X"7f", X"7e", X"7d", X"7f", X"2f", X"2e", X"2d", X"2d", X"2b", X"2a", X"2f", X"2d", X"2f", X"2d", X"2c", X"2b", X"28", X"28", X"2b", X"2c", X"2c", X"2d", X"2a", X"2c", X"29", X"2c", X"2e", X"2f", X"2f", X"2f", X"2d", X"29", X"2e", X"2b", X"2e", X"2d", X"2b", X"2c", X"2a", X"29", X"2c", X"2e", X"2f", X"30", X"2c", X"2b", X"27", X"2b", X"2c", X"2d", X"2f", X"39", X"7f", X"7f", X"7d", X"7d", X"7e", X"7a", X"7c", X"7a", X"79", X"7c", X"7f", X"7f", X"7f", X"7d", X"7f", X"7f", X"7f", X"7f", X"57", X"33", X"2c", X"2f", X"2a", X"2c", X"2d", X"2e", X"2e", X"2a", X"29", X"2c", X"2b", X"2a", X"2d", X"2b", X"2e", X"2b", X"2c", X"2a", X"2c", X"2a", X"2a", X"2d", X"2b", X"2c", X"2d", X"2e", X"2c", X"2d", X"2e", X"2b", X"2b", X"2b", X"2c", X"2b", X"2e", X"2e", X"2e", X"2d", X"31", X"2c", X"34", X"57", X"7f", X"7d", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7d", X"7a", X"7f", X"7f", X"7f", X"7b", X"7f", X"7f", X"7e", X"7d", X"7d", X"7c", X"7b", X"7f", X"7f", X"30", X"31", X"2d", X"2d", X"29", X"2c", X"2c", X"2a", X"2b", X"2b", X"2e", X"2c", X"2a", X"2d", X"2b", X"2e", X"31", X"31", X"32", X"32", X"2f", X"30", X"2c", X"2a", X"2c", X"29", X"2b", X"2a", X"2a", X"2b", X"2a", X"2b", X"2c", X"29", X"29", X"2b", X"2e", X"32", X"7f", X"7f", X"7a", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7a", X"7f", X"7f", X"7f", X"79", X"7a", X"7d", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7c", X"7d", X"7d", X"7f", X"7f", X"54", X"35", X"29", X"2e", X"2c", X"2d", X"2c", X"2a", X"2d", X"2e", X"2e", X"2d", X"2d", X"2b", X"2c", X"2a", X"29", X"2a", X"2b", X"2c", X"2d", X"2d", X"2d", X"2c", X"2b", X"2b", X"2c", X"2b", X"2c", X"28", X"35", X"58", X"7f", X"7f", X"7e", X"7c", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7e", X"7d", X"7d", X"7d", X"7f", X"7e", X"7c", X"7d", X"7c", X"7d", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7d", X"7f", X"7f", X"7d", X"7f", X"7f", X"7b", X"5c", X"49", X"3c", X"2f", X"2a", X"2a", X"27", X"25", X"28", X"28", X"2b", X"2c", X"2d", X"2c", X"2c", X"2a", X"29", X"2a", X"2c", X"2d", X"32", X"3f", X"4c", X"58", X"77", X"7f", X"7f", X"7d", X"7d", X"7d", X"7e", X"7f", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7e", X"7d", X"7c", X"7c", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7b", X"7a", X"7c", X"7e", X"7f", X"7f", X"64", X"5d", X"47", X"36", X"38", X"2f", X"31", X"3a", X"38", X"49", X"5f", X"66", X"7f", X"7f", X"7f", X"7c", X"7c", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7f", X"7d", X"7d", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7d", X"7f", X"7f", X"7d", X"7d", X"7d", X"7d", X"7f", X"7b", X"7e", X"7d", X"7d", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7e", X"7f", X"7f", X"7f", X"7f", X"7f", X"7e", X"7d", X"7d", X"7c", X"7f", X"7f", X"7e", X"7f", X"7d", X"7d", X"7d", X"7d", X"7f", X"7f", X"7f", X"7d", X"7d", X"7c", X"7b", X"7d", X"7f", X"7f", X"7f", X"7d", X"7d", X"7c", X"7e", X"7f", X"7d", X"7e", X"7e", X"7e", X"7f", X"7f"
    );

begin

    RAM_address <= (others => '0');

    re <= '1';

    -- ROM
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (re = '1') then
                R <= std_logic_vector(resize(r_rom(to_integer(unsigned(pixel_y) * 64 + unsigned(pixel_x))), 7));
                G <= std_logic_vector(resize(g_rom(to_integer(unsigned(pixel_y) * 64 + unsigned(pixel_x))), 7));
                B <= std_logic_vector(resize(b_rom(to_integer(unsigned(pixel_y) * 64 + unsigned(pixel_x))), 7));
            end if;
        end if;
    end process;

end Behavioral;

