library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity VGA_pixel_gen is
    Port(clk      : in  STD_LOGIC;
         pixel_x  : in  STD_LOGIC_VECTOR(10 downto 0);
         pixel_y  : in  STD_LOGIC_VECTOR(10 downto 0);
         video_on : in  STD_LOGIC;
         R, G, B  : out STD_LOGIC_VECTOR(6 downto 0));
end VGA_pixel_gen;

architecture Behavioral of VGA_pixel_gen is
    signal R_int, G_int, B_int : STD_LOGIC_VECTOR(7 downto 0) := (others => '0');
    signal re                  : std_logic                    := '1';
    type RomType is array (0 to 4095) of std_logic_vector(7 downto 0);

    constant r_rom : RomType := (
        X"42", X"49", X"34", X"4a", X"7e", X"6b", X"5d", X"5d", X"5e", X"68", X"71", X"70", X"5e", X"4e", X"5e", X"56", X"57", X"52", X"49", X"4d", X"52", X"46", X"2e", X"1e", X"11", X"08", X"00", X"07", X"1e", X"00", X"04", X"04", X"14", X"00", X"00", X"11", X"09", X"00", X"00", X"0a", X"04", X"00", X"00", X"02", X"05", X"04", X"00", X"2c", X"0c", X"65", X"6d", X"70", X"6e", X"6b", X"68", X"64", X"63", X"5e", X"5b", X"5b", X"54", X"52", X"6a", X"6b", X"6a", X"3d", X"0b", X"29", X"63", X"53", X"6f", X"76", X"54", X"57", X"5c", X"57", X"58", X"47", X"5b", X"58", X"55", X"50", X"57", X"4f", X"4a", X"34", X"1d", X"15", X"10", X"09", X"07", X"04", X"03", X"06", X"00", X"03", X"16", X"05", X"10", X"00", X"01", X"04", X"07", X"03", X"00", X"00", X"02", X"00", X"0a", X"17", X"00", X"00", X"00", X"05", X"13", X"61", X"63", X"69", X"68", X"66", X"61", X"5e", X"5b", X"56", X"55", X"65", X"6c", X"6f", X"69", X"3e", X"1e", X"18", X"30", X"60", X"68", X"70", X"6d", X"74", X"64", X"66", X"5a", X"4c", X"39", X"5a", X"56", X"52", X"52", X"4e", X"42", X"36", X"2a", X"19", X"14", X"0e", X"0c", X"0c", X"2b", X"15", X"11", X"14", X"04", X"1e", X"13", X"09", X"0a", X"03", X"03", X"0a", X"04", X"03", X"0b", X"07", X"00", X"04", X"01", X"02", X"02", X"03", X"03", X"01", X"07", X"0b", X"0c", X"23", X"36", X"3b", X"38", X"2d", X"23", X"2d", X"3e", X"3b", X"4d", X"41", X"48", X"46", X"32", X"34", X"75", X"5c", X"57", X"79", X"57", X"62", X"62", X"5c", X"54", X"4c", X"45", X"4f", X"59", X"48", X"44", X"2c", X"29", X"22", X"17", X"13", X"11", X"10", X"14", X"16", X"1a", X"19", X"04", X"07", X"1c", X"00", X"1b", X"0d", X"07", X"0a", X"00", X"13", X"01", X"0b", X"08", X"06", X"04", X"04", X"04", X"01", X"01", X"04", X"07", X"0a", X"0b", X"0b", X"09", X"03", X"29", X"41", X"4c", X"68", X"6c", X"6a", X"4f", X"45", X"59", X"49", X"3f", X"38", X"29", X"61", X"67", X"59", X"51", X"49", X"5c", X"5d", X"5b", X"5e", X"69", X"5f", X"40", X"47", X"3f", X"33", X"29", X"29", X"1b", X"20", X"21", X"49", X"1b", X"1a", X"21", X"13", X"1b", X"10", X"00", X"15", X"0a", X"06", X"04", X"0b", X"00", X"03", X"09", X"08", X"05", X"00", X"03", X"03", X"01", X"08", X"05", X"05", X"07", X"03", X"38", X"56", X"5c", X"5f", X"57", X"56", X"56", X"6e", X"6b", X"6f", X"31", X"3f", X"47", X"49", X"45", X"55", X"43", X"47", X"57", X"67", X"6b", X"6e", X"6f", X"60", X"76", X"74", X"68", X"4c", X"57", X"45", X"41", X"3b", X"37", X"35", X"33", X"35", X"46", X"35", X"20", X"1d", X"1e", X"23", X"1a", X"00", X"18", X"09", X"02", X"03", X"04", X"06", X"09", X"00", X"0b", X"02", X"00", X"00", X"02", X"02", X"00", X"00", X"04", X"04", X"58", X"65", X"6c", X"6c", X"67", X"63", X"5d", X"5a", X"57", X"68", X"6a", X"6d", X"10", X"0d", X"11", X"06", X"24", X"41", X"2a", X"2d", X"66", X"51", X"69", X"68", X"55", X"71", X"72", X"6c", X"56", X"3f", X"50", X"46", X"45", X"46", X"41", X"4a", X"44", X"4d", X"55", X"2b", X"25", X"21", X"1c", X"1b", X"11", X"00", X"20", X"0b", X"08", X"05", X"0f", X"09", X"03", X"00", X"0a", X"04", X"07", X"04", X"02", X"00", X"00", X"01", X"07", X"0b", X"3b", X"67", X"6a", X"6a", X"65", X"63", X"63", X"5a", X"58", X"5d", X"6a", X"6d", X"65", X"71", X"45", X"30", X"46", X"26", X"13", X"25", X"56", X"5a", X"56", X"5f", X"53", X"6e", X"6f", X"69", X"61", X"46", X"5e", X"4f", X"44", X"53", X"57", X"54", X"59", X"5a", X"53", X"3e", X"1e", X"32", X"26", X"44", X"19", X"04", X"00", X"24", X"17", X"00", X"00", X"19", X"08", X"00", X"0f", X"04", X"01", X"00", X"00", X"01", X"04", X"05", X"03", X"05", X"05", X"0c", X"12", X"5d", X"62", X"63", X"5d", X"5b", X"55", X"55", X"6b", X"6e", X"68", X"78", X"53", X"5e", X"2d", X"12", X"04", X"32", X"54", X"73", X"65", X"75", X"47", X"66", X"66", X"5c", X"58", X"4d", X"3f", X"3a", X"3b", X"50", X"68", X"66", X"5f", X"5a", X"4a", X"48", X"3e", X"3f", X"51", X"27", X"1a", X"10", X"17", X"0c", X"13", X"13", X"19", X"09", X"02", X"00", X"0f", X"05", X"04", X"04", X"03", X"02", X"01", X"01", X"00", X"00", X"00", X"00", X"01", X"14", X"1c", X"43", X"5b", X"61", X"59", X"55", X"5d", X"6b", X"6c", X"58", X"61", X"60", X"26", X"0f", X"10", X"2d", X"5c", X"61", X"71", X"58", X"50", X"48", X"52", X"63", X"4b", X"51", X"4d", X"4b", X"52", X"5f", X"6b", X"66", X"45", X"47", X"53", X"4a", X"52", X"4f", X"4f", X"2d", X"28", X"22", X"37", X"34", X"22", X"09", X"1d", X"04", X"03", X"00", X"00", X"13", X"0a", X"01", X"01", X"01", X"03", X"00", X"04", X"04", X"4e", X"6c", X"74", X"6e", X"5e", X"41", X"3a", X"4c", X"59", X"5c", X"57", X"5b", X"54", X"56", X"70", X"5b", X"5c", X"13", X"1f", X"22", X"6a", X"60", X"5e", X"63", X"55", X"73", X"6b", X"6b", X"6c", X"4e", X"5c", X"5c", X"55", X"65", X"72", X"62", X"63", X"5d", X"6a", X"5a", X"66", X"6b", X"60", X"48", X"39", X"35", X"44", X"23", X"27", X"0e", X"00", X"17", X"0b", X"01", X"01", X"05", X"07", X"0a", X"0f", X"12", X"0d", X"02", X"09", X"68", X"71", X"76", X"77", X"79", X"76", X"6c", X"65", X"60", X"40", X"54", X"57", X"51", X"64", X"50", X"5e", X"5b", X"35", X"2a", X"28", X"2c", X"27", X"40", X"61", X"5f", X"71", X"6b", X"74", X"74", X"67", X"4f", X"4b", X"49", X"60", X"61", X"52", X"6a", X"53", X"50", X"5f", X"4f", X"53", X"52", X"60", X"61", X"5e", X"4f", X"53", X"55", X"58", X"2b", X"2d", X"1e", X"00", X"23", X"14", X"0c", X"05", X"00", X"0b", X"0a", X"05", X"03", X"66", X"74", X"78", X"79", X"78", X"77", X"79", X"79", X"76", X"70", X"63", X"4c", X"62", X"5f", X"6a", X"65", X"66", X"5c", X"48", X"35", X"36", X"1d", X"1f", X"3e", X"7a", X"6c", X"72", X"61", X"72", X"76", X"7f", X"5a", X"53", X"57", X"6a", X"69", X"5f", X"60", X"75", X"5d", X"4c", X"37", X"6b", X"50", X"4a", X"5a", X"5f", X"5c", X"6b", X"5b", X"46", X"32", X"22", X"00", X"1b", X"09", X"09", X"00", X"00", X"16", X"0b", X"05", X"03", X"03", X"72", X"70", X"7f", X"7f", X"7a", X"7b", X"7f", X"7b", X"7a", X"77", X"6e", X"67", X"6d", X"6c", X"67", X"5e", X"61", X"5c", X"57", X"3d", X"56", X"3a", X"15", X"2e", X"5e", X"4a", X"7f", X"64", X"63", X"7f", X"6b", X"65", X"63", X"79", X"6a", X"5f", X"55", X"28", X"35", X"2a", X"2e", X"1e", X"2b", X"4a", X"69", X"61", X"51", X"5c", X"3b", X"38", X"45", X"44", X"37", X"15", X"12", X"06", X"08", X"00", X"10", X"0a", X"05", X"01", X"01", X"00", X"61", X"76", X"7a", X"79", X"7e", X"7c", X"7e", X"7f", X"79", X"74", X"71", X"55", X"7a", X"7f", X"5a", X"63", X"54", X"51", X"47", X"4e", X"3f", X"4a", X"28", X"2a", X"14", X"1d", X"4b", X"4e", X"7f", X"71", X"6f", X"56", X"53", X"67", X"69", X"52", X"42", X"37", X"46", X"2e", X"2a", X"33", X"4a", X"41", X"54", X"5f", X"4e", X"52", X"3c", X"3d", X"46", X"58", X"24", X"12", X"0e", X"04", X"03", X"02", X"16", X"0c", X"03", X"01", X"05", X"11", X"0c", X"6f", X"74", X"79", X"77", X"78", X"76", X"75", X"73", X"66", X"5f", X"63", X"69", X"6b", X"53", X"4c", X"4f", X"53", X"5d", X"45", X"3c", X"4a", X"5d", X"39", X"28", X"1c", X"27", X"69", X"4d", X"65", X"64", X"7d", X"57", X"60", X"47", X"38", X"3a", X"48", X"3c", X"50", X"51", X"41", X"3e", X"2b", X"25", X"19", X"21", X"2b", X"2a", X"3f", X"61", X"5b", X"46", X"48", X"20", X"19", X"0d", X"06", X"00", X"15", X"11", X"09", X"17", X"06", X"04", X"06", X"6f", X"76", X"78", X"78", X"79", X"6b", X"3b", X"31", X"59", X"5e", X"62", X"5c", X"2f", X"33", X"48", X"42", X"73", X"4d", X"52", X"38", X"32", X"3e", X"4f", X"4b", X"17", X"1d", X"32", X"42", X"6d", X"78", X"4d", X"48", X"30", X"25", X"3d", X"3e", X"43", X"3f", X"44", X"51", X"4e", X"41", X"35", X"3b", X"0e", X"24", X"31", X"55", X"6c", X"49", X"54", X"26", X"27", X"19", X"00", X"14", X"0b", X"00", X"00", X"1e", X"09", X"07", X"02", X"00", X"06", X"06", X"04", X"0d", X"22", X"14", X"5b", X"65", X"63", X"5b", X"56", X"68", X"1d", X"28", X"4d", X"52", X"35", X"29", X"22", X"41", X"33", X"45", X"3a", X"3e", X"1d", X"1f", X"13", X"0f", X"4b", X"2b", X"57", X"18", X"26", X"2e", X"61", X"38", X"29", X"2d", X"15", X"29", X"0b", X"20", X"48", X"3b", X"44", X"34", X"32", X"49", X"58", X"41", X"39", X"49", X"39", X"1f", X"00", X"1f", X"20", X"00", X"18", X"00", X"1b", X"04", X"09", X"05", X"00", X"10", X"0e", X"08", X"59", X"67", X"63", X"5f", X"57", X"4e", X"71", X"73", X"24", X"22", X"2e", X"47", X"53", X"5c", X"49", X"32", X"0d", X"24", X"17", X"0f", X"2e", X"18", X"0c", X"1b", X"08", X"11", X"03", X"08", X"1c", X"31", X"42", X"27", X"0f", X"18", X"1c", X"09", X"07", X"33", X"2d", X"37", X"3d", X"3d", X"43", X"2e", X"36", X"4e", X"47", X"68", X"37", X"22", X"16", X"0a", X"0f", X"1b", X"17", X"01", X"00", X"0d", X"09", X"07", X"01", X"02", X"59", X"64", X"66", X"66", X"60", X"57", X"54", X"74", X"78", X"77", X"28", X"00", X"31", X"31", X"4b", X"5c", X"40", X"18", X"1d", X"16", X"1a", X"1f", X"53", X"35", X"3b", X"19", X"11", X"19", X"0e", X"2f", X"25", X"37", X"61", X"2e", X"1b", X"00", X"0e", X"00", X"43", X"38", X"17", X"2b", X"3a", X"64", X"4a", X"45", X"53", X"4e", X"4c", X"47", X"49", X"2c", X"36", X"38", X"26", X"0a", X"00", X"1e", X"00", X"18", X"10", X"0f", X"0d", X"4d", X"65", X"6a", X"68", X"61", X"5a", X"58", X"7a", X"7c", X"7d", X"7e", X"21", X"00", X"14", X"33", X"64", X"4c", X"3a", X"2d", X"63", X"59", X"62", X"5a", X"45", X"25", X"2f", X"3d", X"41", X"3e", X"44", X"51", X"48", X"56", X"4d", X"27", X"1a", X"32", X"35", X"4a", X"73", X"52", X"19", X"15", X"0e", X"2a", X"3e", X"31", X"62", X"5a", X"5b", X"69", X"43", X"50", X"55", X"48", X"4c", X"4c", X"1a", X"24", X"08", X"16", X"09", X"0f", X"12", X"63", X"69", X"6b", X"65", X"5f", X"5b", X"54", X"77", X"7f", X"7e", X"7c", X"10", X"01", X"20", X"14", X"33", X"40", X"52", X"3f", X"65", X"4f", X"61", X"73", X"71", X"3d", X"43", X"3d", X"4e", X"4c", X"38", X"3a", X"4c", X"42", X"37", X"32", X"4d", X"6e", X"5c", X"60", X"5d", X"54", X"67", X"41", X"33", X"0b", X"2f", X"48", X"4f", X"4e", X"50", X"64", X"63", X"60", X"60", X"57", X"5b", X"5d", X"46", X"40", X"21", X"11", X"1b", X"10", X"0e", X"5e", X"6b", X"6b", X"67", X"5f", X"5a", X"55", X"78", X"7f", X"7f", X"7d", X"1f", X"00", X"1b", X"16", X"3b", X"3c", X"2b", X"3b", X"55", X"4e", X"58", X"58", X"4f", X"3e", X"44", X"31", X"23", X"26", X"30", X"40", X"1b", X"3e", X"3c", X"4a", X"6f", X"64", X"57", X"7b", X"75", X"69", X"68", X"4d", X"37", X"28", X"2f", X"3d", X"40", X"62", X"5c", X"63", X"58", X"5b", X"5e", X"37", X"43", X"46", X"54", X"46", X"30", X"18", X"18", X"09", X"0e", X"03", X"61", X"6b", X"6a", X"6a", X"5b", X"56", X"76", X"78", X"77", X"7a", X"0b", X"1a", X"09", X"10", X"1e", X"3e", X"47", X"53", X"4d", X"53", X"65", X"51", X"5a", X"5a", X"3f", X"38", X"4f", X"4d", X"3d", X"33", X"3d", X"52", X"67", X"5b", X"6a", X"5b", X"59", X"73", X"7a", X"68", X"61", X"4b", X"43", X"37", X"18", X"21", X"35", X"65", X"49", X"61", X"68", X"6a", X"4a", X"27", X"1b", X"2e", X"2c", X"37", X"29", X"12", X"20", X"0f", X"09", X"0c", X"0e", X"60", X"68", X"63", X"63", X"5a", X"65", X"79", X"7e", X"7f", X"08", X"06", X"00", X"2d", X"20", X"3a", X"31", X"43", X"57", X"2d", X"39", X"62", X"52", X"53", X"69", X"51", X"6d", X"4e", X"5d", X"6e", X"6c", X"5e", X"59", X"6c", X"5f", X"4c", X"4c", X"50", X"6b", X"68", X"52", X"7a", X"69", X"29", X"1f", X"21", X"2f", X"44", X"3c", X"59", X"5a", X"4b", X"38", X"2a", X"5f", X"45", X"53", X"45", X"20", X"06", X"15", X"09", X"06", X"00", X"01", X"1e", X"14", X"5a", X"61", X"60", X"57", X"72", X"7a", X"7e", X"0c", X"0e", X"0b", X"07", X"1c", X"00", X"00", X"1c", X"1e", X"15", X"43", X"40", X"33", X"49", X"62", X"4d", X"56", X"5c", X"5d", X"68", X"67", X"5e", X"70", X"68", X"5b", X"62", X"62", X"51", X"68", X"71", X"5f", X"5d", X"44", X"35", X"2e", X"30", X"40", X"03", X"1a", X"16", X"1c", X"10", X"25", X"3e", X"5d", X"44", X"36", X"18", X"0d", X"15", X"0b", X"04", X"05", X"44", X"70", X"6f", X"67", X"40", X"4f", X"62", X"62", X"5a", X"7c", X"7d", X"05", X"03", X"07", X"0c", X"00", X"1c", X"22", X"00", X"0e", X"32", X"00", X"21", X"2e", X"4d", X"4e", X"68", X"4e", X"5e", X"48", X"50", X"4e", X"5b", X"67", X"60", X"5d", X"5f", X"64", X"58", X"73", X"6f", X"78", X"6c", X"6e", X"2f", X"4a", X"3d", X"20", X"16", X"0f", X"13", X"19", X"23", X"45", X"43", X"54", X"51", X"14", X"25", X"13", X"03", X"12", X"06", X"70", X"7a", X"7a", X"7d", X"7f", X"75", X"6d", X"3f", X"6c", X"6b", X"5c", X"72", X"01", X"05", X"02", X"03", X"00", X"18", X"10", X"00", X"06", X"14", X"00", X"17", X"27", X"21", X"29", X"4d", X"34", X"3a", X"40", X"63", X"60", X"4d", X"42", X"40", X"47", X"56", X"60", X"65", X"5c", X"5a", X"5f", X"53", X"53", X"47", X"38", X"26", X"3f", X"3b", X"3f", X"4c", X"4a", X"41", X"3f", X"4d", X"36", X"36", X"25", X"01", X"06", X"0f", X"08", X"00", X"63", X"73", X"76", X"79", X"77", X"77", X"74", X"73", X"78", X"75", X"71", X"5b", X"07", X"04", X"04", X"05", X"21", X"00", X"23", X"00", X"00", X"17", X"0b", X"13", X"0a", X"0e", X"1a", X"21", X"27", X"26", X"46", X"51", X"58", X"47", X"45", X"44", X"51", X"45", X"5d", X"6f", X"70", X"54", X"59", X"5b", X"79", X"58", X"30", X"26", X"47", X"4e", X"37", X"2d", X"1d", X"2b", X"69", X"43", X"42", X"33", X"18", X"10", X"0c", X"0e", X"08", X"05", X"65", X"78", X"77", X"74", X"72", X"6c", X"67", X"68", X"6a", X"6b", X"6d", X"7a", X"6d", X"0b", X"06", X"00", X"07", X"08", X"09", X"16", X"00", X"00", X"11", X"14", X"1f", X"00", X"08", X"1d", X"1e", X"1d", X"40", X"54", X"42", X"3c", X"37", X"41", X"52", X"4f", X"6e", X"74", X"74", X"67", X"62", X"5b", X"54", X"5e", X"40", X"36", X"31", X"40", X"40", X"31", X"24", X"3a", X"5e", X"44", X"37", X"2e", X"2a", X"1e", X"11", X"06", X"05", X"21", X"0a", X"67", X"6f", X"6e", X"69", X"5d", X"3f", X"4c", X"52", X"55", X"53", X"58", X"65", X"07", X"0a", X"0c", X"0a", X"04", X"02", X"05", X"00", X"12", X"10", X"02", X"0f", X"18", X"0e", X"23", X"1f", X"1f", X"21", X"30", X"24", X"2c", X"27", X"3c", X"4d", X"5f", X"6a", X"73", X"6b", X"60", X"79", X"78", X"71", X"5c", X"56", X"2c", X"3e", X"57", X"46", X"57", X"50", X"42", X"49", X"3a", X"38", X"3a", X"1f", X"05", X"13", X"03", X"0b", X"00", X"05", X"03", X"0d", X"27", X"1d", X"48", X"54", X"53", X"72", X"72", X"71", X"70", X"65", X"09", X"0a", X"08", X"08", X"04", X"08", X"00", X"03", X"04", X"00", X"10", X"10", X"00", X"13", X"11", X"09", X"0e", X"3d", X"1e", X"1c", X"25", X"33", X"34", X"46", X"40", X"5b", X"5b", X"5c", X"50", X"50", X"5a", X"6a", X"6a", X"44", X"46", X"3a", X"40", X"19", X"3c", X"29", X"2a", X"52", X"31", X"3c", X"22", X"21", X"0a", X"00", X"1a", X"08", X"06", X"07", X"07", X"40", X"58", X"58", X"58", X"5a", X"73", X"74", X"70", X"70", X"6b", X"52", X"17", X"13", X"05", X"01", X"01", X"00", X"10", X"00", X"00", X"15", X"07", X"17", X"04", X"0a", X"1b", X"28", X"00", X"06", X"11", X"14", X"1b", X"25", X"26", X"41", X"47", X"5f", X"46", X"45", X"50", X"57", X"64", X"5a", X"6a", X"4e", X"3f", X"25", X"38", X"2c", X"45", X"64", X"6a", X"5b", X"4f", X"3f", X"2a", X"00", X"16", X"00", X"13", X"05", X"04", X"07", X"0f", X"10", X"49", X"54", X"54", X"6e", X"71", X"6f", X"6f", X"6e", X"69", X"00", X"1c", X"03", X"00", X"00", X"02", X"00", X"01", X"00", X"1c", X"02", X"00", X"00", X"0a", X"03", X"06", X"0c", X"19", X"00", X"0e", X"15", X"1e", X"26", X"30", X"41", X"49", X"50", X"5c", X"39", X"4b", X"59", X"51", X"5c", X"5c", X"51", X"6a", X"34", X"29", X"2f", X"5f", X"47", X"57", X"5b", X"50", X"2e", X"00", X"2d", X"18", X"08", X"00", X"0d", X"02", X"00", X"01", X"02", X"1b", X"19", X"3e", X"5f", X"6e", X"71", X"70", X"70", X"6e", X"10", X"00", X"24", X"18", X"05", X"02", X"05", X"04", X"19", X"00", X"15", X"1d", X"00", X"02", X"00", X"00", X"00", X"14", X"00", X"10", X"14", X"1b", X"2f", X"43", X"4f", X"53", X"54", X"59", X"3b", X"58", X"63", X"60", X"6d", X"66", X"57", X"2b", X"32", X"47", X"45", X"52", X"52", X"42", X"59", X"2a", X"0b", X"2b", X"13", X"04", X"06", X"00", X"03", X"0c", X"1e", X"51", X"5c", X"5c", X"59", X"56", X"63", X"58", X"70", X"6d", X"68", X"65", X"63", X"65", X"67", X"69", X"64", X"16", X"06", X"01", X"02", X"05", X"05", X"02", X"14", X"00", X"00", X"04", X"0e", X"17", X"07", X"21", X"41", X"4d", X"56", X"47", X"53", X"54", X"57", X"3d", X"4a", X"61", X"71", X"73", X"5d", X"6a", X"3e", X"2f", X"46", X"5b", X"43", X"5f", X"5f", X"5e", X"5a", X"46", X"29", X"0b", X"08", X"00", X"00", X"16", X"06", X"03", X"08", X"4d", X"5e", X"5f", X"5a", X"54", X"6d", X"73", X"6d", X"6c", X"67", X"64", X"5c", X"61", X"67", X"68", X"6c", X"61", X"06", X"00", X"00", X"00", X"04", X"09", X"12", X"0e", X"02", X"15", X"03", X"0a", X"15", X"19", X"1d", X"27", X"2b", X"33", X"46", X"4d", X"62", X"68", X"72", X"6a", X"51", X"6c", X"65", X"5d", X"3b", X"20", X"1a", X"3d", X"4d", X"4e", X"48", X"5c", X"3c", X"30", X"27", X"17", X"04", X"07", X"0d", X"15", X"08", X"04", X"03", X"59", X"60", X"64", X"5a", X"51", X"54", X"5e", X"6c", X"70", X"6f", X"68", X"5d", X"61", X"65", X"64", X"63", X"5a", X"01", X"06", X"06", X"06", X"00", X"03", X"0c", X"09", X"00", X"09", X"0a", X"17", X"19", X"1a", X"1b", X"1c", X"20", X"1c", X"2f", X"43", X"55", X"49", X"5e", X"6b", X"65", X"56", X"6a", X"76", X"2e", X"18", X"59", X"5d", X"50", X"60", X"5e", X"48", X"48", X"1e", X"26", X"15", X"00", X"0c", X"00", X"14", X"0b", X"01", X"0a", X"0b", X"60", X"5f", X"53", X"39", X"4b", X"4c", X"69", X"6c", X"66", X"64", X"52", X"5c", X"5d", X"64", X"64", X"5a", X"06", X"02", X"02", X"03", X"00", X"0a", X"16", X"00", X"00", X"08", X"1b", X"00", X"12", X"1e", X"22", X"25", X"20", X"2c", X"2e", X"40", X"4c", X"39", X"58", X"55", X"54", X"4a", X"29", X"26", X"23", X"2a", X"5c", X"58", X"5f", X"57", X"58", X"63", X"5b", X"57", X"2c", X"12", X"16", X"11", X"09", X"00", X"14", X"06", X"01", X"02", X"00", X"1b", X"11", X"53", X"60", X"67", X"64", X"64", X"6d", X"79", X"51", X"59", X"63", X"63", X"61", X"1b", X"15", X"02", X"02", X"04", X"05", X"0f", X"00", X"0c", X"0a", X"14", X"14", X"15", X"15", X"15", X"17", X"1b", X"25", X"1d", X"35", X"46", X"58", X"46", X"57", X"5b", X"66", X"35", X"48", X"37", X"2a", X"50", X"69", X"77", X"6b", X"62", X"45", X"5a", X"53", X"30", X"25", X"15", X"15", X"00", X"07", X"23", X"12", X"00", X"05", X"0a", X"12", X"00", X"65", X"74", X"7a", X"7f", X"78", X"6c", X"58", X"5f", X"49", X"50", X"56", X"2d", X"09", X"05", X"06", X"03", X"18", X"08", X"08", X"08", X"00", X"0a", X"09", X"08", X"0d", X"1d", X"00", X"13", X"18", X"1d", X"32", X"46", X"45", X"58", X"68", X"70", X"6c", X"48", X"58", X"4b", X"41", X"3a", X"29", X"76", X"63", X"5a", X"52", X"5e", X"4a", X"47", X"46", X"44", X"2d", X"28", X"22", X"1f", X"09", X"37", X"0f", X"00", X"12", X"0c", X"0c", X"61", X"73", X"7e", X"70", X"66", X"58", X"68", X"6c", X"6d", X"32", X"14", X"15", X"11", X"07", X"01", X"00", X"02", X"0b", X"00", X"01", X"0d", X"04", X"01", X"00", X"04", X"09", X"16", X"29", X"01", X"1a", X"33", X"49", X"5b", X"5a", X"59", X"5b", X"4b", X"5e", X"4f", X"4b", X"40", X"47", X"37", X"4b", X"5c", X"55", X"5e", X"6a", X"4f", X"55", X"5f", X"5c", X"4a", X"48", X"44", X"55", X"2a", X"2a", X"26", X"06", X"18", X"06", X"07", X"11", X"47", X"74", X"7f", X"7f", X"7d", X"7e", X"7d", X"6a", X"5f", X"51", X"5a", X"5e", X"53", X"0c", X"08", X"04", X"02", X"04", X"0a", X"02", X"03", X"00", X"0b", X"05", X"04", X"09", X"03", X"25", X"00", X"06", X"18", X"26", X"3a", X"4b", X"58", X"5b", X"4c", X"60", X"65", X"57", X"48", X"59", X"34", X"0e", X"3b", X"78", X"72", X"6c", X"6d", X"5e", X"6f", X"6a", X"55", X"50", X"5e", X"5a", X"51", X"66", X"47", X"3a", X"25", X"07", X"0c", X"08", X"05", X"0b", X"4b", X"60", X"63", X"56", X"4f", X"58", X"60", X"5a", X"5c", X"43", X"13", X"10", X"08", X"03", X"01", X"00", X"06", X"1a", X"00", X"0d", X"00", X"0d", X"02", X"07", X"13", X"00", X"02", X"0b", X"1c", X"24", X"3e", X"4a", X"4e", X"42", X"51", X"60", X"50", X"61", X"44", X"41", X"39", X"36", X"27", X"41", X"50", X"55", X"62", X"60", X"5a", X"6c", X"66", X"62", X"4d", X"4d", X"4e", X"2f", X"42", X"43", X"55", X"2f", X"0f", X"1d", X"12", X"07", X"51", X"50", X"4a", X"6b", X"76", X"78", X"76", X"24", X"08", X"01", X"01", X"01", X"01", X"02", X"04", X"07", X"0c", X"15", X"00", X"02", X"15", X"0c", X"07", X"16", X"00", X"0b", X"14", X"17", X"1c", X"25", X"44", X"4d", X"53", X"65", X"5b", X"51", X"58", X"58", X"61", X"52", X"2e", X"3b", X"47", X"29", X"4a", X"76", X"6c", X"5a", X"65", X"67", X"63", X"50", X"65", X"3c", X"38", X"3f", X"41", X"39", X"2b", X"2d", X"1f", X"10", X"11", X"61", X"6b", X"62", X"69", X"78", X"75", X"7a", X"7c", X"6e", X"71", X"72", X"67", X"05", X"05", X"05", X"02", X"02", X"09", X"15", X"00", X"00", X"0f", X"00", X"20", X"15", X"30", X"1a", X"33", X"31", X"2c", X"36", X"43", X"4b", X"64", X"70", X"61", X"6f", X"6a", X"52", X"36", X"1e", X"1e", X"3d", X"50", X"28", X"1f", X"1e", X"23", X"54", X"59", X"5f", X"72", X"4d", X"37", X"26", X"27", X"3e", X"2b", X"3d", X"42", X"46", X"14", X"1f", X"06", X"46", X"60", X"44", X"47", X"70", X"79", X"7f", X"7b", X"74", X"75", X"74", X"6e", X"43", X"0c", X"1c", X"0b", X"00", X"00", X"00", X"04", X"07", X"12", X"17", X"12", X"1e", X"1f", X"25", X"41", X"58", X"3f", X"46", X"4d", X"59", X"46", X"53", X"4f", X"52", X"41", X"2a", X"18", X"33", X"3a", X"56", X"60", X"3e", X"4c", X"49", X"38", X"38", X"36", X"55", X"53", X"3e", X"23", X"2c", X"61", X"53", X"59", X"53", X"3f", X"47", X"3f", X"2d", X"00", X"0b", X"0c", X"54", X"56", X"73", X"7c", X"76", X"79", X"7e", X"7a", X"77", X"71", X"6d", X"0b", X"0e", X"01", X"11", X"14", X"00", X"10", X"07", X"17", X"00", X"12", X"1f", X"27", X"2d", X"45", X"50", X"5a", X"42", X"54", X"43", X"52", X"52", X"65", X"78", X"3a", X"45", X"48", X"56", X"5e", X"30", X"34", X"33", X"2d", X"27", X"23", X"13", X"1e", X"16", X"0d", X"20", X"2b", X"35", X"4a", X"57", X"52", X"60", X"47", X"4a", X"58", X"30", X"19", X"22", X"0a", X"64", X"6c", X"65", X"58", X"6a", X"6e", X"78", X"7e", X"7e", X"75", X"3a", X"04", X"03", X"03", X"00", X"13", X"19", X"06", X"11", X"0d", X"13", X"1d", X"4a", X"2d", X"3c", X"45", X"59", X"4a", X"66", X"62", X"5b", X"51", X"51", X"6a", X"70", X"3d", X"55", X"5e", X"43", X"3f", X"41", X"46", X"1b", X"27", X"16", X"14", X"25", X"41", X"3d", X"39", X"28", X"39", X"4c", X"49", X"5b", X"48", X"48", X"46", X"68", X"51", X"3d", X"34", X"17", X"12", X"60", X"5d", X"65", X"5f", X"5c", X"5e", X"1b", X"07", X"0d", X"06", X"01", X"07", X"08", X"06", X"05", X"09", X"0f", X"12", X"00", X"23", X"3f", X"40", X"49", X"59", X"50", X"56", X"58", X"5d", X"63", X"71", X"60", X"71", X"5d", X"59", X"4e", X"35", X"2d", X"1f", X"21", X"33", X"21", X"48", X"23", X"4e", X"4c", X"5f", X"4e", X"52", X"4e", X"48", X"5b", X"39", X"58", X"38", X"23", X"43", X"37", X"3c", X"43", X"32", X"36", X"42", X"2f", X"2f", X"65", X"55", X"66", X"6b", X"6b", X"6b", X"54", X"0f", X"17", X"03", X"07", X"03", X"07", X"0e", X"08", X"12", X"26", X"00", X"14", X"28", X"2a", X"57", X"54", X"62", X"51", X"66", X"61", X"59", X"69", X"59", X"5a", X"66", X"55", X"66", X"25", X"1b", X"26", X"26", X"13", X"14", X"40", X"2c", X"29", X"5f", X"70", X"69", X"51", X"52", X"5c", X"54", X"46", X"54", X"19", X"1b", X"2e", X"13", X"28", X"3a", X"3d", X"2b", X"24", X"1b", X"11", X"22", X"61", X"69", X"6c", X"6a", X"67", X"5f", X"68", X"5a", X"0a", X"16", X"05", X"07", X"0b", X"21", X"00", X"17", X"22", X"1c", X"3d", X"54", X"57", X"3e", X"35", X"39", X"65", X"58", X"63", X"62", X"71", X"66", X"43", X"24", X"25", X"22", X"23", X"2a", X"39", X"52", X"4c", X"5f", X"37", X"22", X"1f", X"3c", X"4e", X"5e", X"57", X"5d", X"4a", X"30", X"2c", X"1b", X"33", X"00", X"00", X"1d", X"10", X"00", X"0d", X"22", X"09", X"0e", X"33", X"65", X"64", X"54", X"67", X"69", X"62", X"5d", X"70", X"65", X"10", X"0d", X"17", X"1a", X"3b", X"35", X"20", X"29", X"45", X"30", X"3d", X"62", X"63", X"61", X"5b", X"2e", X"22", X"36", X"3b", X"42", X"31", X"2f", X"3c", X"43", X"3a", X"3d", X"4e", X"3f", X"6f", X"4d", X"4a", X"51", X"3a", X"2f", X"11", X"36", X"5b", X"42", X"3f", X"2a", X"21", X"00", X"29", X"04", X"04", X"06", X"0a", X"05", X"00", X"13", X"00", X"19", X"2a", X"4f", X"43", X"47", X"64", X"6d", X"6a", X"6b", X"62", X"58", X"4f", X"13", X"0e", X"17", X"28", X"3f", X"48", X"45", X"50", X"55", X"58", X"59", X"4e", X"5b", X"53", X"3d", X"2e", X"33", X"4b", X"3c", X"47", X"3e", X"50", X"68", X"35", X"2e", X"20", X"37", X"48", X"52", X"58", X"5f", X"5e", X"5c", X"69", X"2e", X"43", X"51", X"45", X"59", X"4d", X"1f", X"2a", X"07", X"16", X"00", X"13", X"02", X"00", X"22", X"00", X"2a", X"64", X"6a", X"3b", X"3e", X"69", X"77", X"72", X"67", X"6c", X"65", X"62", X"57", X"00", X"12", X"16", X"07", X"14", X"33", X"41", X"40", X"55", X"5f", X"72", X"54", X"51", X"4f", X"45", X"3a", X"24", X"2d", X"35", X"71", X"67", X"5f", X"5f", X"69", X"63", X"70", X"37", X"46", X"51", X"54", X"54", X"50", X"4b", X"4e", X"5e", X"57", X"54", X"55", X"2d", X"25", X"41", X"1d", X"0e", X"0e", X"0b", X"0b", X"09", X"10", X"3e", X"5c", X"59", X"38", X"7b", X"7d", X"6a", X"4d", X"6a", X"79", X"7a", X"76", X"74", X"65", X"5f", X"52", X"67", X"0e", X"14", X"23", X"1a", X"35", X"2a", X"27", X"3f", X"49", X"47", X"6e", X"5a", X"7f", X"4d", X"3f", X"2c", X"5f", X"5d", X"61", X"4b", X"54", X"5f", X"5f", X"72", X"59", X"61", X"59", X"4f", X"54", X"54", X"41", X"2b", X"36", X"2e", X"5a", X"55", X"55", X"44", X"31", X"12", X"33", X"1c", X"00", X"00", X"07", X"15", X"09", X"1e", X"52", X"56", X"5b", X"70", X"70", X"7e", X"5b", X"69", X"74", X"77", X"7d", X"75", X"6b", X"65", X"57", X"70", X"0e", X"10", X"15", X"1a", X"28", X"49", X"34", X"19", X"30", X"24", X"34", X"28", X"18", X"2d", X"40", X"3b", X"42", X"58", X"6f", X"69", X"71", X"57", X"49", X"57", X"5b", X"59", X"4f", X"55", X"2e", X"27", X"1b", X"14", X"26", X"20", X"15", X"44", X"3e", X"41", X"34", X"09", X"01", X"17", X"07", X"21", X"4e", X"10", X"45", X"32", X"4d", X"4d", X"50", X"5d", X"7f", X"4d", X"7b", X"60", X"6a", X"70", X"76", X"75", X"78", X"63", X"56", X"00", X"0d", X"14", X"00", X"23", X"1f", X"41", X"44", X"5c", X"43", X"32", X"11", X"23", X"33", X"28", X"47", X"55", X"60", X"4d", X"54", X"4a", X"4d", X"41", X"5e", X"47", X"30", X"34", X"3b", X"24", X"2b", X"24", X"00", X"2e", X"00", X"00", X"2b", X"08", X"15", X"3e", X"2d", X"2c", X"0e", X"13", X"01", X"6b", X"7b", X"64", X"3a", X"52", X"49", X"5f", X"5e", X"5a", X"6a", X"6a", X"5c", X"5a", X"7c", X"64", X"6c", X"72", X"7f", X"75", X"67", X"03", X"11", X"0f", X"0c", X"20", X"45", X"5c", X"59", X"63", X"39", X"40", X"4c", X"47", X"43", X"5a", X"52", X"49", X"51", X"5d", X"4c", X"4e", X"4c", X"3c", X"54", X"47", X"2c", X"29", X"2f", X"0f", X"05", X"0e", X"12", X"1b", X"0a", X"05", X"00", X"00", X"1c", X"00", X"0a", X"0f", X"0a", X"06", X"18", X"62", X"7c", X"75", X"69", X"5d", X"65", X"6b", X"6e", X"6a", X"5e", X"7f", X"54", X"58", X"59", X"57", X"69", X"72", X"6b", X"7b", X"69", X"00", X"12", X"05", X"0d", X"35", X"59", X"5a", X"6a", X"4a", X"37", X"2d", X"38", X"46", X"3b", X"24", X"36", X"54", X"51", X"6a", X"5c", X"51", X"3b", X"36", X"3f", X"25", X"29", X"20", X"15", X"00", X"15", X"15", X"00", X"14", X"0a", X"00", X"09", X"00", X"00", X"02", X"13", X"09", X"00", X"53", X"2d", X"33", X"60", X"78", X"71", X"5f", X"63", X"65", X"65", X"64", X"61", X"55", X"53", X"52", X"53", X"51", X"57", X"5c", X"65", X"71", X"75", X"02", X"23", X"1d", X"27", X"40", X"30", X"34", X"34", X"2c", X"28", X"54", X"3e", X"48", X"2b", X"2f", X"3d", X"63", X"5b", X"64", X"63", X"58", X"36", X"27", X"15", X"32", X"0b", X"0d", X"16", X"21", X"10", X"05", X"00", X"04", X"10", X"06", X"04", X"05", X"00", X"01", X"14", X"16", X"5a", X"65", X"65", X"5d", X"4f", X"5e", X"73", X"68", X"60", X"66", X"65", X"5d", X"55", X"4e", X"7f", X"75", X"7d", X"7b", X"79", X"73", X"5f", X"61", X"6f", X"12", X"0d", X"12", X"23", X"49", X"2c", X"1c", X"1b", X"31", X"1e", X"23", X"1e", X"49", X"3d", X"36", X"61", X"50", X"58", X"3b", X"5a", X"44", X"2f", X"1d", X"07", X"00", X"2a", X"17", X"16", X"00", X"13", X"00", X"22", X"1e", X"00", X"02", X"02", X"00", X"55", X"5c", X"13", X"2b", X"55", X"59", X"5e", X"59", X"58", X"5e", X"6e", X"7f", X"5b", X"65", X"64", X"5e", X"59", X"6f", X"75", X"78", X"7c", X"7b", X"76", X"7a", X"74", X"6c", X"67", X"14", X"1f", X"30", X"3d", X"35", X"43", X"54", X"45", X"63", X"58", X"40", X"4b", X"2b", X"35", X"41", X"54", X"60", X"58", X"3f", X"5c", X"5a", X"3d", X"1c", X"0a", X"1b", X"0b", X"0a", X"09", X"17", X"00", X"00", X"15", X"0b", X"04", X"01", X"11", X"65", X"69", X"7d", X"74", X"2d", X"57", X"5b", X"58", X"57", X"76", X"77", X"6f", X"5b", X"7f", X"5f", X"59", X"55", X"5a", X"71", X"78", X"78", X"75", X"7e", X"7e", X"7e", X"7b", X"76", X"73", X"40", X"40", X"53", X"40", X"34", X"45", X"66", X"59", X"5d", X"70", X"62", X"65", X"3d", X"3e", X"31", X"4e", X"64", X"6b", X"62", X"52", X"49", X"29", X"23", X"0e", X"00", X"1d", X"09", X"06", X"12", X"00", X"00", X"0e", X"04", X"0b", X"06", X"04", X"62", X"77", X"7b", X"7f", X"74", X"69", X"5c", X"4f", X"7a", X"7b", X"7a", X"76", X"71", X"69", X"58", X"7f", X"54", X"68", X"6d", X"73", X"77", X"7d", X"7a", X"7c", X"7c", X"7a", X"76", X"74"
    );

    constant g_rom : RomType := (
        X"17", X"27", X"21", X"3e", X"71", X"4c", X"1b", X"0b", X"0b", X"0d", X"06", X"04", X"00", X"01", X"27", X"2b", X"2e", X"2c", X"24", X"2a", X"2f", X"25", X"10", X"09", X"09", X"0a", X"08", X"24", X"5a", X"4b", X"60", X"57", X"4a", X"1a", X"1c", X"34", X"2c", X"2a", X"3d", X"56", X"54", X"51", X"4e", X"49", X"3e", X"38", X"31", X"53", X"1c", X"65", X"63", X"60", X"5b", X"58", X"52", X"4e", X"49", X"41", X"38", X"34", X"2a", X"21", X"2f", X"2b", X"36", X"22", X"21", X"47", X"5e", X"34", X"3c", X"37", X"0e", X"0c", X"0c", X"06", X"05", X"01", X"29", X"32", X"2d", X"29", X"2f", X"27", X"1f", X"12", X"0c", X"10", X"0f", X"0c", X"0a", X"07", X"02", X"06", X"08", X"0c", X"19", X"18", X"47", X"46", X"42", X"3b", X"32", X"28", X"24", X"27", X"2f", X"31", X"4e", X"5e", X"3c", X"35", X"2e", X"28", X"23", X"65", X"5b", X"59", X"53", X"4e", X"47", X"42", X"3c", X"31", X"27", X"2f", X"2e", X"2c", X"37", X"1e", X"20", X"34", X"5e", X"7a", X"49", X"2c", X"15", X"13", X"05", X"09", X"02", X"01", X"00", X"2c", X"30", X"2c", X"28", X"20", X"11", X"0c", X"11", X"0e", X"0d", X"0d", X"0e", X"0c", X"1e", X"07", X"0d", X"1d", X"20", X"4d", X"56", X"51", X"49", X"3e", X"3e", X"4a", X"4e", X"58", X"6a", X"65", X"42", X"4c", X"4b", X"4b", X"41", X"3d", X"3d", X"35", X"2e", X"27", X"1d", X"2b", X"37", X"3a", X"37", X"2f", X"27", X"32", X"40", X"3c", X"1f", X"10", X"10", X"1c", X"27", X"30", X"60", X"31", X"13", X"26", X"00", X"07", X"02", X"00", X"00", X"00", X"00", X"08", X"0d", X"04", X"15", X"0b", X"0e", X"10", X"0f", X"10", X"0d", X"0c", X"0e", X"11", X"18", X"1b", X"08", X"0c", X"1f", X"14", X"53", X"5d", X"61", X"66", X"52", X"63", X"4b", X"57", X"59", X"5a", X"57", X"59", X"5b", X"5c", X"5e", X"63", X"67", X"6e", X"74", X"6c", X"57", X"37", X"3e", X"38", X"26", X"31", X"30", X"2c", X"38", X"33", X"51", X"42", X"2d", X"34", X"48", X"74", X"3e", X"12", X"08", X"00", X"0c", X"0a", X"04", X"01", X"03", X"03", X"06", X"1f", X"17", X"0f", X"05", X"0e", X"0f", X"14", X"07", X"30", X"14", X"1b", X"20", X"11", X"19", X"1f", X"1d", X"5f", X"6a", X"73", X"77", X"73", X"46", X"46", X"55", X"61", X"68", X"69", X"6e", X"71", X"72", X"79", X"71", X"64", X"50", X"34", X"4c", X"55", X"49", X"44", X"3b", X"31", X"20", X"2f", X"2a", X"2b", X"1d", X"26", X"1f", X"18", X"0d", X"20", X"1b", X"29", X"40", X"40", X"1e", X"10", X"10", X"00", X"05", X"03", X"03", X"00", X"21", X"1e", X"1b", X"15", X"0e", X"0c", X"0c", X"10", X"22", X"1a", X"17", X"1c", X"19", X"1f", X"16", X"13", X"65", X"77", X"79", X"7b", X"70", X"60", X"4b", X"30", X"69", X"70", X"70", X"75", X"79", X"77", X"6e", X"5f", X"4a", X"30", X"66", X"5f", X"59", X"52", X"4c", X"45", X"3a", X"31", X"25", X"2e", X"2c", X"2c", X"4b", X"49", X"4e", X"2d", X"1e", X"2f", X"2b", X"2c", X"51", X"20", X"17", X"06", X"00", X"0d", X"05", X"02", X"01", X"00", X"24", X"23", X"1d", X"19", X"0b", X"13", X"10", X"21", X"32", X"15", X"1d", X"22", X"1d", X"1c", X"10", X"11", X"6d", X"75", X"78", X"6e", X"63", X"4f", X"3f", X"3a", X"6f", X"7a", X"7b", X"76", X"70", X"64", X"57", X"4a", X"3f", X"2f", X"46", X"62", X"59", X"55", X"4f", X"49", X"42", X"34", X"2e", X"2c", X"2f", X"2c", X"55", X"72", X"68", X"5b", X"5c", X"36", X"2a", X"2e", X"3d", X"28", X"11", X"0d", X"00", X"0c", X"03", X"01", X"08", X"00", X"27", X"21", X"16", X"1e", X"14", X"11", X"21", X"2b", X"25", X"16", X"01", X"1a", X"10", X"32", X"10", X"0f", X"1a", X"66", X"61", X"42", X"25", X"41", X"35", X"35", X"75", X"79", X"75", X"70", X"70", X"71", X"71", X"71", X"70", X"6d", X"61", X"4f", X"2f", X"60", X"55", X"4e", X"45", X"3e", X"30", X"24", X"2e", X"2b", X"3f", X"56", X"40", X"59", X"35", X"2b", X"30", X"50", X"41", X"42", X"29", X"2f", X"00", X"11", X"06", X"00", X"00", X"00", X"01", X"02", X"00", X"03", X"06", X"09", X"23", X"2f", X"1c", X"1d", X"16", X"1a", X"2a", X"0b", X"10", X"0f", X"14", X"09", X"11", X"26", X"52", X"4f", X"3f", X"35", X"6e", X"75", X"79", X"7c", X"79", X"75", X"6f", X"6a", X"62", X"5c", X"54", X"51", X"56", X"5f", X"52", X"5d", X"4f", X"43", X"39", X"2d", X"25", X"2b", X"27", X"1b", X"33", X"4d", X"39", X"37", X"39", X"47", X"55", X"3d", X"31", X"0d", X"07", X"00", X"04", X"15", X"00", X"07", X"03", X"00", X"00", X"04", X"03", X"05", X"00", X"07", X"08", X"00", X"15", X"1d", X"24", X"0c", X"13", X"11", X"24", X"23", X"1b", X"1b", X"59", X"53", X"4c", X"40", X"35", X"57", X"6c", X"72", X"6e", X"65", X"5a", X"48", X"3c", X"29", X"5f", X"6c", X"69", X"66", X"65", X"53", X"52", X"59", X"49", X"3a", X"2b", X"2c", X"03", X"0b", X"2c", X"34", X"63", X"2e", X"31", X"27", X"5a", X"3a", X"20", X"1a", X"0f", X"27", X"0f", X"0d", X"14", X"00", X"02", X"00", X"00", X"07", X"0c", X"00", X"00", X"00", X"0f", X"03", X"14", X"21", X"22", X"12", X"08", X"0d", X"27", X"11", X"1c", X"18", X"19", X"57", X"59", X"55", X"4f", X"51", X"54", X"5a", X"62", X"62", X"52", X"36", X"26", X"75", X"75", X"71", X"6b", X"6a", X"67", X"60", X"62", X"61", X"3e", X"4b", X"42", X"36", X"13", X"02", X"11", X"25", X"2a", X"3a", X"40", X"42", X"33", X"39", X"40", X"2b", X"2f", X"19", X"11", X"0e", X"11", X"02", X"03", X"00", X"11", X"0e", X"00", X"14", X"00", X"08", X"2e", X"22", X"16", X"08", X"06", X"08", X"14", X"0f", X"1a", X"21", X"2b", X"09", X"1b", X"22", X"15", X"5b", X"70", X"71", X"54", X"39", X"53", X"4e", X"3c", X"2c", X"7c", X"7d", X"78", X"75", X"75", X"73", X"71", X"6f", X"69", X"68", X"68", X"4e", X"53", X"47", X"05", X"05", X"10", X"1a", X"25", X"25", X"2d", X"27", X"44", X"5b", X"6b", X"43", X"3e", X"1c", X"17", X"15", X"2a", X"0a", X"06", X"08", X"13", X"12", X"10", X"19", X"31", X"2a", X"36", X"28", X"47", X"1a", X"04", X"09", X"08", X"09", X"26", X"23", X"19", X"16", X"1a", X"1b", X"71", X"74", X"67", X"50", X"36", X"5c", X"52", X"47", X"3a", X"28", X"7c", X"6b", X"79", X"7e", X"7b", X"7c", X"7a", X"74", X"74", X"75", X"70", X"68", X"69", X"65", X"08", X"00", X"07", X"17", X"33", X"24", X"32", X"25", X"28", X"4b", X"62", X"38", X"59", X"2f", X"24", X"36", X"19", X"11", X"11", X"2c", X"20", X"2d", X"4d", X"3a", X"51", X"44", X"39", X"22", X"2e", X"3b", X"35", X"1a", X"0c", X"26", X"21", X"24", X"1d", X"18", X"18", X"1d", X"5c", X"66", X"54", X"40", X"60", X"5d", X"56", X"4a", X"3a", X"27", X"74", X"7d", X"7c", X"78", X"7c", X"79", X"78", X"7c", X"7d", X"7d", X"7c", X"5d", X"79", X"7b", X"2f", X"2c", X"05", X"0a", X"28", X"3d", X"22", X"33", X"27", X"41", X"42", X"45", X"49", X"34", X"5d", X"41", X"35", X"18", X"15", X"2f", X"40", X"3c", X"45", X"3f", X"40", X"1e", X"10", X"17", X"37", X"32", X"42", X"4e", X"3d", X"48", X"3e", X"33", X"1a", X"27", X"0b", X"0b", X"14", X"17", X"22", X"34", X"5d", X"5f", X"5a", X"50", X"40", X"39", X"23", X"79", X"77", X"77", X"76", X"74", X"70", X"6f", X"72", X"6a", X"66", X"67", X"63", X"60", X"22", X"12", X"01", X"10", X"42", X"36", X"19", X"20", X"35", X"1f", X"26", X"2d", X"44", X"7a", X"37", X"3e", X"42", X"5b", X"30", X"47", X"50", X"41", X"1f", X"22", X"22", X"3a", X"35", X"25", X"24", X"26", X"47", X"4b", X"50", X"48", X"26", X"1a", X"19", X"0e", X"11", X"29", X"13", X"1a", X"18", X"22", X"2e", X"5b", X"5c", X"55", X"5e", X"42", X"30", X"20", X"78", X"73", X"6e", X"6a", X"68", X"65", X"4c", X"44", X"58", X"4e", X"45", X"3a", X"0f", X"0b", X"10", X"0c", X"50", X"34", X"3b", X"27", X"2a", X"3a", X"43", X"49", X"2f", X"3c", X"42", X"47", X"67", X"6e", X"48", X"47", X"34", X"24", X"29", X"19", X"10", X"07", X"0e", X"1e", X"18", X"1c", X"34", X"54", X"39", X"41", X"1e", X"24", X"2b", X"08", X"25", X"08", X"19", X"20", X"14", X"3e", X"37", X"35", X"3b", X"65", X"53", X"53", X"49", X"3f", X"38", X"33", X"34", X"44", X"62", X"43", X"5a", X"49", X"42", X"34", X"2a", X"3a", X"1b", X"1c", X"2f", X"32", X"23", X"1e", X"16", X"2e", X"14", X"20", X"13", X"27", X"27", X"3c", X"35", X"31", X"65", X"41", X"6b", X"29", X"35", X"2d", X"3e", X"16", X"23", X"40", X"3b", X"4e", X"1c", X"1a", X"27", X"0f", X"18", X"14", X"29", X"43", X"3f", X"1b", X"08", X"19", X"17", X"13", X"0c", X"46", X"48", X"2b", X"66", X"53", X"6a", X"54", X"62", X"65", X"65", X"70", X"5d", X"3b", X"5f", X"54", X"49", X"40", X"34", X"23", X"3b", X"38", X"18", X"0d", X"08", X"18", X"1f", X"34", X"3a", X"39", X"25", X"49", X"42", X"2f", X"30", X"21", X"41", X"66", X"53", X"5c", X"4f", X"3e", X"25", X"21", X"2a", X"1e", X"2c", X"51", X"63", X"55", X"50", X"63", X"2e", X"24", X"2b", X"27", X"23", X"10", X"23", X"32", X"0c", X"2b", X"16", X"14", X"13", X"11", X"1e", X"45", X"6c", X"69", X"4c", X"6f", X"77", X"74", X"5d", X"42", X"6b", X"5c", X"56", X"50", X"45", X"33", X"21", X"39", X"3a", X"39", X"63", X"19", X"28", X"0b", X"15", X"2b", X"22", X"1b", X"4b", X"53", X"4a", X"34", X"3f", X"14", X"23", X"13", X"25", X"41", X"43", X"53", X"1a", X"16", X"41", X"26", X"40", X"3a", X"50", X"3e", X"79", X"5e", X"27", X"25", X"1e", X"3d", X"22", X"20", X"36", X"27", X"09", X"00", X"11", X"01", X"13", X"22", X"1e", X"14", X"1a", X"4f", X"36", X"69", X"65", X"58", X"3d", X"65", X"65", X"5c", X"54", X"48", X"3a", X"2e", X"3f", X"3a", X"3b", X"3d", X"6b", X"2d", X"21", X"1e", X"33", X"1e", X"2d", X"2f", X"60", X"4c", X"45", X"40", X"45", X"2a", X"27", X"29", X"22", X"1a", X"1f", X"27", X"11", X"24", X"32", X"26", X"36", X"53", X"3f", X"4b", X"76", X"6a", X"58", X"53", X"25", X"2c", X"3c", X"23", X"3c", X"1c", X"01", X"10", X"03", X"18", X"18", X"08", X"0c", X"21", X"16", X"3e", X"31", X"4e", X"4b", X"49", X"2e", X"68", X"5d", X"57", X"52", X"47", X"39", X"28", X"3e", X"40", X"3d", X"3a", X"4a", X"33", X"42", X"17", X"0c", X"11", X"3f", X"2f", X"43", X"1a", X"18", X"34", X"57", X"31", X"2a", X"1d", X"26", X"28", X"23", X"29", X"34", X"33", X"40", X"3f", X"4b", X"5c", X"38", X"37", X"39", X"41", X"6f", X"5f", X"62", X"2b", X"21", X"29", X"37", X"2c", X"0e", X"0f", X"07", X"03", X"06", X"0d", X"2b", X"35", X"14", X"18", X"19", X"2a", X"55", X"4d", X"30", X"6a", X"65", X"5b", X"54", X"46", X"3a", X"2a", X"3d", X"3f", X"40", X"3e", X"4d", X"27", X"3a", X"20", X"25", X"21", X"22", X"2b", X"25", X"09", X"08", X"16", X"35", X"2d", X"20", X"1d", X"43", X"4b", X"2d", X"32", X"20", X"4d", X"4e", X"48", X"42", X"23", X"19", X"3f", X"39", X"3f", X"5e", X"5d", X"5d", X"47", X"2e", X"2d", X"32", X"44", X"17", X"10", X"0c", X"1f", X"39", X"1d", X"29", X"29", X"33", X"2c", X"28", X"2d", X"53", X"50", X"46", X"25", X"64", X"5d", X"52", X"4e", X"3a", X"2d", X"42", X"3f", X"3c", X"3e", X"69", X"6a", X"39", X"23", X"16", X"24", X"29", X"26", X"05", X"03", X"1a", X"08", X"0e", X"1c", X"1e", X"2c", X"51", X"59", X"50", X"40", X"35", X"33", X"2f", X"14", X"1c", X"0c", X"0d", X"2b", X"37", X"2c", X"2c", X"34", X"5d", X"5b", X"1c", X"21", X"4d", X"70", X"22", X"21", X"28", X"38", X"31", X"2b", X"3c", X"51", X"32", X"2c", X"1a", X"1e", X"67", X"73", X"6c", X"59", X"31", X"66", X"5f", X"4d", X"46", X"35", X"35", X"3f", X"3a", X"38", X"79", X"70", X"5b", X"68", X"23", X"1b", X"06", X"14", X"2c", X"04", X"10", X"2e", X"08", X"0b", X"3c", X"2b", X"3a", X"11", X"18", X"2a", X"35", X"23", X"08", X"15", X"10", X"03", X"06", X"09", X"1b", X"1d", X"1a", X"5e", X"72", X"3d", X"21", X"2a", X"58", X"69", X"3a", X"43", X"45", X"3e", X"3b", X"27", X"44", X"18", X"1e", X"1e", X"20", X"2b", X"5e", X"64", X"5f", X"5a", X"5f", X"6b", X"39", X"62", X"52", X"42", X"2e", X"42", X"41", X"41", X"67", X"62", X"50", X"41", X"4a", X"1a", X"0c", X"20", X"1b", X"09", X"2d", X"1b", X"00", X"0f", X"2e", X"14", X"09", X"03", X"02", X"0b", X"08", X"00", X"0e", X"07", X"00", X"0b", X"11", X"00", X"0b", X"16", X"15", X"2e", X"3b", X"36", X"1d", X"2b", X"67", X"3d", X"50", X"49", X"4d", X"35", X"33", X"32", X"31", X"12", X"14", X"18", X"3f", X"60", X"58", X"45", X"2f", X"5b", X"79", X"75", X"72", X"4a", X"4e", X"54", X"42", X"2a", X"3f", X"39", X"5b", X"58", X"5c", X"60", X"50", X"68", X"5b", X"20", X"3a", X"51", X"06", X"18", X"1d", X"2f", X"1d", X"2b", X"0c", X"17", X"00", X"04", X"00", X"05", X"07", X"00", X"00", X"03", X"09", X"00", X"0f", X"12", X"2b", X"3a", X"61", X"2d", X"3b", X"2b", X"14", X"1c", X"32", X"38", X"24", X"1a", X"2d", X"1f", X"27", X"33", X"1c", X"47", X"44", X"3e", X"4d", X"34", X"7f", X"7c", X"7b", X"7b", X"7c", X"76", X"76", X"43", X"5d", X"4c", X"2f", X"3d", X"3a", X"46", X"53", X"5b", X"4e", X"60", X"43", X"2a", X"4c", X"54", X"19", X"21", X"24", X"14", X"10", X"2d", X"0b", X"0b", X"0d", X"2b", X"23", X"0f", X"05", X"00", X"00", X"04", X"09", X"0f", X"0e", X"0d", X"0f", X"13", X"36", X"43", X"41", X"2f", X"3b", X"29", X"1b", X"20", X"1b", X"1e", X"32", X"40", X"0b", X"0f", X"22", X"18", X"30", X"43", X"3d", X"2b", X"75", X"78", X"77", X"75", X"72", X"75", X"78", X"7a", X"7c", X"71", X"5e", X"40", X"2c", X"34", X"4b", X"53", X"68", X"3a", X"50", X"25", X"3c", X"4b", X"18", X"0f", X"09", X"0b", X"10", X"15", X"1d", X"15", X"24", X"23", X"21", X"11", X"1b", X"1b", X"1f", X"03", X"04", X"0b", X"0f", X"00", X"05", X"12", X"3d", X"3a", X"41", X"35", X"23", X"20", X"26", X"30", X"2a", X"2c", X"47", X"11", X"11", X"10", X"10", X"23", X"39", X"4a", X"43", X"31", X"70", X"71", X"6b", X"67", X"66", X"62", X"5e", X"5e", X"5c", X"5e", X"67", X"76", X"79", X"28", X"42", X"50", X"68", X"71", X"76", X"73", X"36", X"2a", X"65", X"71", X"6b", X"1c", X"18", X"1c", X"1e", X"13", X"21", X"2a", X"16", X"10", X"0c", X"11", X"18", X"02", X"07", X"02", X"05", X"00", X"0b", X"10", X"13", X"37", X"47", X"42", X"1a", X"1d", X"28", X"28", X"2c", X"42", X"4d", X"25", X"13", X"24", X"5b", X"6f", X"67", X"58", X"47", X"4f", X"1e", X"69", X"65", X"60", X"5a", X"53", X"3e", X"46", X"39", X"31", X"2e", X"33", X"76", X"25", X"44", X"5e", X"70", X"77", X"79", X"71", X"3b", X"5e", X"77", X"71", X"74", X"5e", X"20", X"1a", X"12", X"0e", X"0d", X"1a", X"0f", X"13", X"08", X"0d", X"03", X"01", X"00", X"06", X"05", X"00", X"0d", X"11", X"19", X"26", X"53", X"38", X"2f", X"33", X"0f", X"1b", X"21", X"1e", X"2e", X"1e", X"0e", X"19", X"21", X"22", X"43", X"47", X"5e", X"57", X"54", X"4c", X"50", X"5b", X"38", X"48", X"35", X"21", X"37", X"31", X"2d", X"2b", X"71", X"2b", X"55", X"6d", X"77", X"73", X"69", X"54", X"62", X"68", X"63", X"72", X"5e", X"33", X"21", X"0e", X"07", X"09", X"30", X"11", X"12", X"14", X"0c", X"02", X"13", X"03", X"09", X"00", X"06", X"00", X"02", X"10", X"22", X"38", X"3a", X"42", X"1a", X"22", X"1b", X"44", X"1d", X"1d", X"54", X"31", X"27", X"1b", X"4a", X"4c", X"32", X"6d", X"76", X"79", X"69", X"4a", X"54", X"4e", X"41", X"33", X"26", X"35", X"32", X"2c", X"2e", X"29", X"71", X"47", X"66", X"69", X"64", X"5d", X"4e", X"55", X"39", X"42", X"6f", X"5b", X"48", X"2b", X"3b", X"49", X"49", X"09", X"0b", X"0e", X"11", X"14", X"19", X"0a", X"0c", X"08", X"24", X"08", X"00", X"04", X"0b", X"19", X"0d", X"33", X"43", X"46", X"23", X"34", X"2d", X"3d", X"43", X"31", X"0d", X"07", X"17", X"23", X"18", X"4a", X"39", X"71", X"71", X"71", X"67", X"55", X"30", X"49", X"3b", X"28", X"37", X"33", X"30", X"2f", X"2c", X"26", X"45", X"69", X"54", X"48", X"45", X"49", X"4e", X"56", X"4b", X"71", X"4a", X"39", X"2c", X"3d", X"45", X"4e", X"4e", X"48", X"0b", X"0b", X"13", X"15", X"12", X"12", X"1d", X"22", X"26", X"2c", X"00", X"04", X"0d", X"04", X"0e", X"1e", X"34", X"62", X"32", X"25", X"20", X"3d", X"07", X"08", X"0a", X"0e", X"0d", X"07", X"63", X"63", X"4c", X"42", X"6b", X"65", X"57", X"47", X"2e", X"38", X"30", X"40", X"3b", X"34", X"2e", X"27", X"26", X"24", X"51", X"2c", X"3f", X"2d", X"25", X"2e", X"3d", X"42", X"57", X"3a", X"51", X"53", X"24", X"2e", X"3b", X"47", X"4b", X"4e", X"0c", X"10", X"11", X"0f", X"14", X"20", X"28", X"2d", X"2f", X"2f", X"00", X"0e", X"0f", X"0b", X"22", X"35", X"50", X"30", X"23", X"31", X"30", X"31", X"17", X"02", X"28", X"12", X"15", X"5a", X"6b", X"68", X"58", X"42", X"44", X"41", X"3f", X"5d", X"4f", X"3f", X"31", X"2a", X"38", X"28", X"32", X"2b", X"29", X"28", X"4c", X"50", X"52", X"5a", X"5c", X"22", X"2e", X"3c", X"46", X"51", X"57", X"53", X"5c", X"2e", X"38", X"3b", X"46", X"3f", X"0d", X"0f", X"1f", X"24", X"28", X"1a", X"2a", X"2c", X"2b", X"08", X"03", X"0c", X"11", X"17", X"12", X"3e", X"42", X"3c", X"34", X"3a", X"22", X"2f", X"10", X"0a", X"19", X"1a", X"11", X"0b", X"1f", X"28", X"2b", X"5b", X"52", X"41", X"21", X"4d", X"51", X"47", X"38", X"27", X"34", X"33", X"2b", X"2b", X"25", X"23", X"41", X"46", X"4d", X"52", X"5c", X"63", X"24", X"35", X"45", X"4e", X"5a", X"5c", X"59", X"48", X"2e", X"32", X"12", X"0f", X"1a", X"1a", X"19", X"1b", X"15", X"11", X"16", X"0b", X"0c", X"04", X"03", X"03", X"00", X"28", X"26", X"35", X"3a", X"33", X"2e", X"46", X"3d", X"28", X"0d", X"21", X"16", X"1a", X"1c", X"1d", X"1d", X"31", X"45", X"56", X"4e", X"3f", X"23", X"62", X"52", X"4b", X"40", X"34", X"33", X"31", X"2f", X"2b", X"28", X"22", X"38", X"40", X"4d", X"53", X"58", X"5e", X"1b", X"33", X"41", X"50", X"58", X"5e", X"5e", X"4b", X"26", X"1f", X"11", X"17", X"17", X"19", X"1d", X"1f", X"20", X"12", X"15", X"1a", X"1f", X"02", X"02", X"0b", X"15", X"1b", X"48", X"70", X"45", X"34", X"62", X"47", X"10", X"0d", X"0b", X"02", X"1b", X"04", X"1a", X"1b", X"11", X"38", X"2d", X"5a", X"54", X"42", X"37", X"21", X"5c", X"55", X"54", X"37", X"3a", X"2a", X"34", X"2c", X"24", X"21", X"34", X"40", X"45", X"51", X"57", X"5f", X"24", X"36", X"45", X"53", X"59", X"61", X"5c", X"2f", X"3e", X"3f", X"44", X"14", X"1b", X"1d", X"1c", X"1f", X"1b", X"20", X"12", X"19", X"20", X"00", X"07", X"06", X"1f", X"39", X"46", X"52", X"3d", X"2c", X"3c", X"1e", X"12", X"01", X"02", X"19", X"26", X"32", X"11", X"10", X"38", X"48", X"40", X"3c", X"5f", X"56", X"4e", X"4f", X"4f", X"5c", X"35", X"5d", X"53", X"50", X"4e", X"50", X"59", X"65", X"31", X"3a", X"45", X"4c", X"58", X"28", X"3e", X"41", X"4d", X"59", X"60", X"61", X"2c", X"34", X"25", X"25", X"18", X"14", X"16", X"17", X"1b", X"1a", X"19", X"07", X"14", X"1d", X"25", X"06", X"09", X"17", X"48", X"24", X"2c", X"1e", X"26", X"45", X"3d", X"32", X"16", X"10", X"09", X"2b", X"27", X"0f", X"16", X"11", X"17", X"11", X"2d", X"5d", X"5d", X"53", X"70", X"72", X"64", X"33", X"70", X"6c", X"71", X"77", X"6a", X"53", X"2c", X"29", X"35", X"41", X"4e", X"34", X"27", X"37", X"49", X"4f", X"61", X"4b", X"41", X"3e", X"32", X"46", X"55", X"59", X"5a", X"54", X"0b", X"0d", X"0e", X"0c", X"13", X"1a", X"0a", X"0b", X"07", X"08", X"0b", X"02", X"3c", X"3e", X"27", X"24", X"28", X"70", X"3a", X"19", X"02", X"0c", X"01", X"04", X"07", X"0f", X"0a", X"10", X"0e", X"1c", X"20", X"60", X"40", X"36", X"6f", X"66", X"43", X"7c", X"79", X"77", X"67", X"52", X"33", X"35", X"2c", X"27", X"3d", X"31", X"5a", X"6f", X"6d", X"6e", X"6a", X"6b", X"69", X"54", X"5f", X"72", X"70", X"70", X"69", X"6b", X"69", X"61", X"4f", X"0a", X"0c", X"17", X"22", X"2f", X"2d", X"27", X"20", X"06", X"0c", X"0b", X"2f", X"31", X"28", X"23", X"5c", X"67", X"2f", X"1c", X"20", X"00", X"02", X"0b", X"0a", X"00", X"0b", X"13", X"2c", X"0a", X"10", X"20", X"20", X"49", X"48", X"4a", X"45", X"65", X"75", X"75", X"7b", X"76", X"74", X"69", X"45", X"31", X"3a", X"45", X"4b", X"58", X"3a", X"57", X"6d", X"76", X"7a", X"74", X"55", X"52", X"57", X"74", X"7a", X"78", X"70", X"59", X"66", X"15", X"12", X"0d", X"09", X"14", X"25", X"2d", X"27", X"09", X"0c", X"17", X"2a", X"28", X"32", X"20", X"28", X"56", X"67", X"41", X"22", X"14", X"00", X"0c", X"09", X"00", X"00", X"09", X"04", X"03", X"25", X"16", X"17", X"19", X"1a", X"3d", X"53", X"50", X"3b", X"62", X"5f", X"52", X"3e", X"30", X"36", X"3b", X"40", X"4d", X"4d", X"38", X"53", X"5f", X"64", X"6b", X"71", X"71", X"6f", X"38", X"4d", X"35", X"71", X"77", X"7c", X"6f", X"1e", X"09", X"0e", X"14", X"09", X"14", X"12", X"0d", X"00", X"07", X"0f", X"0c", X"40", X"35", X"35", X"2e", X"27", X"22", X"4c", X"4d", X"1f", X"12", X"0c", X"02", X"10", X"0b", X"0a", X"08", X"27", X"3c", X"20", X"2b", X"16", X"2d", X"28", X"31", X"6d", X"68", X"39", X"66", X"4c", X"2f", X"3e", X"3c", X"36", X"32", X"58", X"40", X"40", X"4b", X"59", X"66", X"71", X"79", X"79", X"76", X"6d", X"38", X"4d", X"50", X"28", X"17", X"2d", X"0d", X"06", X"09", X"12", X"10", X"04", X"11", X"0b", X"05", X"0a", X"00", X"00", X"18", X"31", X"4f", X"4f", X"28", X"18", X"2b", X"33", X"58", X"61", X"3c", X"16", X"15", X"11", X"16", X"18", X"3d", X"21", X"24", X"2a", X"37", X"44", X"34", X"21", X"1d", X"37", X"3b", X"67", X"57", X"3f", X"3b", X"44", X"3c", X"3b", X"3b", X"56", X"5c", X"62", X"68", X"23", X"3e", X"54", X"62", X"6e", X"70", X"67", X"3d", X"4b", X"50", X"16", X"22", X"0e", X"25", X"0c", X"1f", X"11", X"07", X"12", X"14", X"03", X"0a", X"08", X"00", X"14", X"36", X"5e", X"5d", X"37", X"1f", X"19", X"2c", X"24", X"33", X"3f", X"38", X"40", X"29", X"1e", X"3a", X"37", X"33", X"27", X"36", X"64", X"4a", X"36", X"29", X"2c", X"15", X"54", X"41", X"58", X"5e", X"40", X"35", X"42", X"3e", X"43", X"40", X"6d", X"6d", X"6c", X"6f", X"56", X"32", X"55", X"4b", X"37", X"33", X"38", X"44", X"52", X"55", X"3d", X"23", X"20", X"15", X"0c", X"1f", X"2f", X"14", X"1c", X"1f", X"24", X"06", X"07", X"0e", X"33", X"38", X"2d", X"15", X"17", X"18", X"3b", X"45", X"19", X"29", X"2f", X"32", X"52", X"4f", X"4c", X"4b", X"5c", X"41", X"24", X"3d", X"1b", X"29", X"42", X"30", X"1a", X"22", X"4a", X"3e", X"57", X"46", X"5d", X"39", X"3d", X"3a", X"37", X"3a", X"7a", X"78", X"78", X"77", X"77", X"25", X"41", X"46", X"60", X"63", X"35", X"53", X"57", X"59", X"11", X"16", X"1f", X"1d", X"14", X"21", X"2a", X"2c", X"07", X"10", X"00", X"06", X"00", X"1b", X"4f", X"23", X"2d", X"2e", X"36", X"42", X"20", X"2b", X"29", X"23", X"1b", X"23", X"2a", X"48", X"4c", X"3b", X"34", X"2b", X"26", X"23", X"0d", X"09", X"40", X"2d", X"11", X"21", X"17", X"20", X"4c", X"37", X"74", X"67", X"51", X"35", X"37", X"32", X"71", X"78", X"7b", X"7d", X"55", X"32", X"45", X"52", X"45", X"67", X"69", X"42", X"25", X"0d", X"13", X"14", X"2e", X"03", X"0a", X"11", X"28", X"0d", X"0c", X"00", X"03", X"03", X"0d", X"3a", X"5b", X"2c", X"2d", X"2d", X"13", X"16", X"25", X"37", X"1c", X"3e", X"47", X"3f", X"28", X"30", X"29", X"2c", X"27", X"30", X"24", X"0f", X"1a", X"0d", X"1a", X"22", X"47", X"34", X"28", X"34", X"38", X"3a", X"71", X"5c", X"56", X"42", X"34", X"31", X"50", X"36", X"2e", X"29", X"33", X"45", X"4b", X"4b", X"45", X"55", X"78", X"6d", X"22", X"1e", X"27", X"14", X"09", X"11", X"09", X"0b", X"06", X"01", X"00", X"0b", X"00", X"18", X"12", X"28", X"40", X"32", X"1a", X"1b", X"4a", X"5d", X"1e", X"3a", X"29", X"52", X"37", X"45", X"40", X"43", X"2d", X"22", X"3a", X"15", X"2b", X"0e", X"07", X"2a", X"13", X"1e", X"3a", X"2a", X"18", X"29", X"33", X"36", X"55", X"33", X"34", X"2e", X"26", X"23", X"6b", X"38", X"62", X"59", X"4c", X"41", X"44", X"3d", X"1e", X"20", X"3b", X"12", X"18", X"1a", X"07", X"2d", X"2f", X"32", X"06", X"0d", X"0a", X"04", X"15", X"09", X"0f", X"30", X"41", X"68", X"2f", X"2d", X"3f", X"49", X"41", X"3b", X"49", X"2f", X"39", X"5a", X"37", X"15", X"00", X"0b", X"24", X"27", X"1d", X"34", X"07", X"1a", X"44", X"22", X"12", X"15", X"1a", X"1d", X"3b", X"47", X"41", X"3e", X"51", X"3c", X"30", X"26", X"23", X"1a", X"5c", X"68", X"4a", X"71", X"5e", X"5b", X"55", X"59", X"19", X"20", X"20", X"10", X"24", X"2c", X"1c", X"0b", X"26", X"2f", X"42", X"1e", X"17", X"13", X"31", X"40", X"42", X"36", X"34", X"28", X"17", X"1c", X"38", X"4f", X"37", X"48", X"2b", X"27", X"39", X"43", X"1a", X"0e", X"0a", X"1c", X"18", X"0b", X"0d", X"18", X"5f", X"3c", X"32", X"54", X"41", X"2f", X"41", X"5c", X"4b", X"48", X"55", X"72", X"5b", X"36", X"31", X"27", X"1c", X"16", X"5e", X"69", X"3f", X"45", X"36", X"20", X"28", X"1a", X"0d", X"16", X"26", X"09", X"10", X"28", X"15", X"1e", X"42", X"2e", X"28", X"42", X"48", X"4d", X"36", X"28", X"21", X"22", X"1e", X"20", X"2b", X"1b", X"4c", X"23", X"0b", X"1b", X"28", X"36", X"23", X"3d", X"40", X"19", X"1c", X"14", X"1b", X"13", X"67", X"52", X"46", X"44", X"48", X"4d", X"54", X"70", X"50", X"54", X"41", X"4f", X"3a", X"39", X"51", X"4c", X"30", X"25", X"1d", X"14", X"65", X"36", X"4a", X"47", X"29", X"22", X"1f", X"0f", X"0b", X"08", X"0a", X"0a", X"00", X"1a", X"2c", X"28", X"21", X"25", X"33", X"24", X"39", X"37", X"4b", X"6d", X"47", X"44", X"2d", X"3e", X"49", X"3f", X"1c", X"0d", X"03", X"10", X"41", X"17", X"27", X"31", X"20", X"32", X"26", X"0d", X"40", X"39", X"59", X"4e", X"6c", X"4f", X"2c", X"48", X"2c", X"61", X"7d", X"75", X"47", X"39", X"40", X"3f", X"3c", X"31", X"2f", X"24", X"1c", X"0d", X"4d", X"68", X"6f", X"44", X"14", X"16", X"27", X"26", X"37", X"3c", X"43", X"1a", X"0a", X"15", X"30", X"34", X"16", X"21", X"34", X"66", X"41", X"23", X"11", X"19", X"1e", X"41", X"25", X"2f", X"12", X"03", X"06", X"09", X"0d", X"10", X"11", X"0e", X"1f", X"3d", X"37", X"33", X"32", X"18", X"37", X"53", X"5b", X"64", X"69", X"5c", X"59", X"64", X"6a", X"46", X"7b", X"73", X"5b", X"32", X"3b", X"3f", X"3e", X"3b", X"3d", X"2b", X"1e", X"0d", X"78", X"2f", X"52", X"5a", X"23", X"2e", X"31", X"25", X"1f", X"24", X"33", X"5c", X"3c", X"60", X"24", X"2b", X"43", X"76", X"47", X"2c", X"08", X"05", X"0a", X"02", X"10", X"08", X"36", X"37", X"12", X"13", X"21", X"1b", X"11", X"1d", X"0c", X"2c", X"15", X"1a", X"20", X"29", X"24", X"61", X"67", X"51", X"46", X"4f", X"6c", X"52", X"3b", X"57", X"53", X"54", X"67", X"65", X"6f", X"3f", X"35", X"34", X"37", X"3e", X"3a", X"2d", X"1e", X"0c", X"7c", X"27", X"46", X"45", X"1f", X"17", X"31", X"2d", X"38", X"57", X"34", X"46", X"4f", X"37", X"24", X"2c", X"39", X"30", X"15", X"0e", X"00", X"08", X"02", X"00", X"0f", X"11", X"08", X"09", X"2a", X"15", X"16", X"0f", X"09", X"1e", X"1f", X"0b", X"21", X"17", X"24", X"2d", X"1f", X"2f", X"56", X"43", X"42", X"65", X"2c", X"5d", X"3c", X"48", X"38", X"36", X"48", X"6f", X"32", X"57", X"2f", X"30", X"2f", X"38", X"41", X"45", X"25", X"13", X"2a", X"3f", X"54", X"33", X"3c", X"14", X"0a", X"0c", X"4c", X"42", X"27", X"19", X"58", X"65", X"24", X"2b", X"3f", X"3e", X"0e", X"06", X"00", X"09", X"0b", X"2e", X"15", X"00", X"08", X"17", X"0f", X"21", X"1d", X"06", X"55", X"1a", X"27", X"47", X"12", X"0d", X"22", X"27", X"62", X"63", X"67", X"3f", X"7c", X"7c", X"73", X"47", X"4b", X"30", X"34", X"2e", X"2f", X"3f", X"33", X"25", X"29", X"4a", X"26", X"2b", X"33", X"3f", X"2c", X"1a", X"67", X"6c", X"57", X"37", X"23", X"22", X"12", X"15", X"4d", X"33", X"2a", X"27", X"16", X"13", X"36", X"33", X"27", X"22", X"15", X"03", X"1b", X"21", X"0c", X"29", X"27", X"16", X"1a", X"26", X"0b", X"08", X"1a", X"39", X"6e", X"67", X"4a", X"3d", X"3f", X"6d", X"37", X"4c", X"55", X"55", X"59", X"57", X"74", X"78", X"72", X"5c", X"3d", X"33", X"29", X"25", X"22", X"1d", X"5d", X"23", X"18", X"18", X"1e", X"33", X"39", X"2e", X"3a", X"26", X"66", X"6e", X"41", X"22", X"1a", X"24", X"1e", X"42", X"50", X"4b", X"2a", X"23", X"24", X"1f", X"20", X"30", X"30", X"10", X"0e", X"04", X"1a", X"13", X"09", X"17", X"09", X"17", X"14", X"1f", X"2d", X"54", X"4f", X"2d", X"66", X"5e", X"36", X"46", X"3b", X"44", X"61", X"72", X"4e", X"2d", X"6d", X"3e", X"47", X"71", X"7b", X"65", X"3f", X"32", X"29", X"21", X"1c", X"1a", X"15", X"14", X"0e", X"0d", X"08", X"0c", X"12", X"1d", X"31", X"38", X"3d", X"52", X"33", X"29", X"34", X"1e", X"24", X"2d", X"31", X"28", X"39", X"1b", X"2b", X"21", X"42", X"40", X"2c", X"03", X"04", X"0b", X"14", X"0a", X"11", X"0c", X"2b", X"06", X"0a", X"24", X"4e", X"4f", X"48", X"46", X"4b", X"58", X"4d", X"47", X"3e", X"3d", X"57", X"64", X"42", X"6a", X"5d", X"56", X"59", X"53", X"66", X"71", X"4d", X"31", X"27", X"20", X"19", X"15", X"11", X"43", X"14", X"12", X"10", X"11", X"0f", X"07", X"19", X"30", X"45", X"31", X"16", X"17", X"3b", X"2c", X"37", X"3b", X"3d", X"23", X"2d", X"1e", X"2e", X"1e", X"2a", X"49", X"0e", X"0b", X"00", X"29", X"16", X"0c", X"0c", X"0e", X"0f", X"69", X"71", X"6e", X"28", X"44", X"34", X"5d", X"5e", X"40", X"44", X"3a", X"23", X"6f", X"78", X"31", X"4c", X"6a", X"56", X"4c", X"40", X"3d", X"43", X"54", X"6e", X"3a", X"26", X"18", X"12", X"0a", X"15", X"14", X"11", X"11", X"10", X"0c", X"0f", X"0f", X"11", X"12", X"6c", X"57", X"24", X"1c", X"2d", X"43", X"4b", X"33", X"45", X"40", X"3c", X"4b", X"1f", X"25", X"37", X"38", X"1d", X"08", X"00", X"29", X"2f", X"1d", X"0a", X"10", X"44", X"56", X"72", X"75", X"6b", X"4c", X"42", X"72", X"73", X"68", X"51", X"46", X"77", X"6b", X"7b", X"77", X"3d", X"62", X"4f", X"38", X"27", X"3b", X"37", X"35", X"33", X"5c", X"2f", X"1f", X"12", X"0c", X"12", X"13", X"11", X"0d", X"13", X"11", X"0e", X"0d", X"0c", X"0b", X"1c", X"15", X"1a", X"12", X"27", X"36", X"2f", X"0f", X"11", X"25", X"1b", X"3a", X"48", X"59", X"34", X"30", X"1c", X"0f", X"08", X"05", X"15", X"0b", X"12", X"14", X"10", X"5e", X"64", X"6b", X"6d", X"59", X"51", X"71", X"72", X"74", X"5c", X"3c", X"72", X"70", X"74", X"78", X"70", X"60", X"47", X"29", X"42", X"3a", X"3b", X"37", X"30", X"2d", X"2b", X"56", X"0f", X"16", X"13", X"11", X"0b", X"0f", X"0c", X"0f", X"10", X"10", X"0f", X"0f"
    );

    constant b_rom : RomType := (
        X"1b", X"2e", X"32", X"3c", X"41", X"15", X"05", X"0b", X"1c", X"32", X"45", X"48", X"33", X"31", X"60", X"6c", X"76", X"76", X"6e", X"73", X"7a", X"6c", X"51", X"47", X"4a", X"45", X"39", X"46", X"6c", X"53", X"64", X"5f", X"61", X"38", X"39", X"4e", X"3a", X"27", X"26", X"32", X"31", X"2b", X"27", X"24", X"22", X"22", X"24", X"3e", X"00", X"23", X"0c", X"02", X"03", X"03", X"01", X"01", X"05", X"03", X"00", X"02", X"00", X"00", X"08", X"04", X"34", X"27", X"36", X"4e", X"3b", X"00", X"17", X"1e", X"01", X"07", X"10", X"15", X"27", X"30", X"65", X"74", X"74", X"72", X"7c", X"71", X"5f", X"4d", X"4c", X"51", X"4f", X"4b", X"46", X"3e", X"33", X"33", X"31", X"3c", X"59", X"4e", X"58", X"44", X"3f", X"37", X"2d", X"1f", X"1a", X"1a", X"22", X"25", X"45", X"53", X"2a", X"20", X"18", X"08", X"00", X"1f", X"08", X"02", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"0b", X"05", X"00", X"47", X"33", X"43", X"43", X"36", X"3c", X"17", X"09", X"08", X"16", X"15", X"27", X"30", X"33", X"2d", X"63", X"7c", X"7f", X"77", X"66", X"4b", X"45", X"53", X"55", X"59", X"56", X"4d", X"47", X"5d", X"4b", X"56", X"62", X"57", X"71", X"64", X"59", X"5b", X"51", X"4d", X"54", X"52", X"59", X"6e", X"5f", X"2c", X"2a", X"25", X"23", X"1f", X"1d", X"1d", X"16", X"12", X"0a", X"00", X"08", X"0b", X"09", X"09", X"06", X"07", X"12", X"1b", X"14", X"30", X"24", X"2a", X"35", X"3a", X"2c", X"38", X"00", X"00", X"21", X"16", X"2f", X"36", X"35", X"2f", X"2b", X"27", X"33", X"40", X"38", X"48", X"42", X"52", X"5b", X"5d", X"5c", X"53", X"50", X"53", X"5c", X"6d", X"6c", X"4a", X"49", X"61", X"4a", X"6c", X"66", X"67", X"6c", X"5e", X"6a", X"45", X"42", X"34", X"2f", X"2d", X"2e", X"2f", X"2d", X"2d", X"31", X"33", X"38", X"3d", X"38", X"2c", X"0f", X"15", X"10", X"00", X"09", X"02", X"00", X"2b", X"21", X"36", X"2a", X"28", X"2b", X"25", X"4b", X"22", X"03", X"08", X"0d", X"2c", X"33", X"2d", X"33", X"42", X"44", X"3a", X"4e", X"4c", X"44", X"3a", X"49", X"56", X"5f", X"4c", X"74", X"5e", X"69", X"72", X"65", X"6c", X"63", X"45", X"73", X"73", X"74", X"77", X"77", X"52", X"48", X"3c", X"35", X"36", X"31", X"37", X"39", X"3b", X"42", X"3a", X"32", X"29", X"0b", X"14", X"12", X"03", X"01", X"03", X"02", X"00", X"09", X"03", X"03", X"3d", X"47", X"41", X"33", X"1b", X"26", X"22", X"23", X"21", X"1e", X"10", X"0e", X"14", X"14", X"44", X"4d", X"3c", X"33", X"65", X"65", X"5e", X"51", X"42", X"3e", X"41", X"4a", X"60", X"61", X"6a", X"74", X"72", X"74", X"69", X"50", X"7b", X"77", X"76", X"78", X"73", X"64", X"4d", X"23", X"3d", X"36", X"3a", X"3e", X"3f", X"3b", X"30", X"2b", X"28", X"0a", X"28", X"12", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"03", X"02", X"42", X"44", X"50", X"38", X"36", X"49", X"3f", X"30", X"39", X"06", X"11", X"15", X"19", X"44", X"4c", X"48", X"33", X"2d", X"60", X"65", X"5f", X"57", X"46", X"4e", X"52", X"63", X"73", X"5c", X"72", X"7b", X"75", X"6c", X"54", X"41", X"7f", X"7f", X"7d", X"75", X"70", X"58", X"3d", X"24", X"41", X"3f", X"42", X"3d", X"3b", X"33", X"2d", X"27", X"23", X"09", X"07", X"13", X"08", X"03", X"00", X"00", X"01", X"00", X"00", X"01", X"02", X"00", X"05", X"28", X"2b", X"37", X"5f", X"47", X"33", X"26", X"1c", X"01", X"00", X"0c", X"15", X"3d", X"45", X"3f", X"30", X"1f", X"53", X"54", X"4b", X"55", X"4c", X"4c", X"61", X"6b", X"64", X"58", X"48", X"62", X"56", X"75", X"54", X"48", X"3e", X"7e", X"76", X"57", X"42", X"57", X"39", X"21", X"44", X"3e", X"3d", X"3a", X"3a", X"38", X"36", X"38", X"3b", X"3c", X"33", X"20", X"00", X"24", X"0e", X"05", X"05", X"07", X"02", X"00", X"05", X"01", X"02", X"18", X"03", X"2d", X"2c", X"31", X"31", X"41", X"15", X"0f", X"02", X"1f", X"0a", X"34", X"31", X"26", X"24", X"1e", X"1b", X"1c", X"1e", X"30", X"44", X"50", X"6e", X"74", X"5a", X"57", X"54", X"59", X"67", X"4b", X"5a", X"58", X"52", X"45", X"55", X"5f", X"6c", X"58", X"44", X"29", X"45", X"3b", X"3e", X"41", X"43", X"40", X"3a", X"34", X"2c", X"27", X"24", X"24", X"2b", X"33", X"1f", X"22", X"0b", X"00", X"01", X"00", X"00", X"06", X"0d", X"00", X"01", X"1e", X"22", X"2c", X"34", X"34", X"24", X"07", X"10", X"00", X"05", X"03", X"06", X"16", X"01", X"12", X"20", X"27", X"2b", X"3a", X"49", X"4b", X"33", X"34", X"35", X"30", X"4c", X"57", X"60", X"4c", X"5e", X"60", X"6f", X"6e", X"68", X"56", X"6f", X"55", X"50", X"3d", X"25", X"38", X"3e", X"3b", X"35", X"30", X"2f", X"26", X"23", X"09", X"24", X"1f", X"12", X"0d", X"16", X"0d", X"15", X"21", X"10", X"05", X"00", X"03", X"00", X"00", X"0b", X"0f", X"48", X"20", X"31", X"1d", X"30", X"09", X"01", X"06", X"00", X"1c", X"0a", X"0c", X"17", X"0a", X"2e", X"34", X"24", X"31", X"42", X"33", X"34", X"2b", X"30", X"25", X"45", X"5b", X"5f", X"4e", X"40", X"45", X"67", X"56", X"68", X"56", X"39", X"66", X"64", X"5d", X"55", X"54", X"55", X"57", X"5c", X"57", X"44", X"19", X"00", X"24", X"0f", X"02", X"00", X"02", X"02", X"00", X"08", X"0f", X"00", X"0e", X"0b", X"01", X"2c", X"10", X"0d", X"17", X"1e", X"32", X"40", X"38", X"0f", X"08", X"11", X"01", X"0c", X"04", X"0d", X"11", X"11", X"06", X"11", X"0d", X"10", X"0a", X"01", X"1c", X"05", X"06", X"21", X"13", X"12", X"17", X"34", X"42", X"4b", X"45", X"54", X"5e", X"6c", X"4d", X"62", X"63", X"48", X"7d", X"7f", X"75", X"56", X"32", X"3a", X"2d", X"1b", X"00", X"2c", X"19", X"0b", X"03", X"04", X"02", X"03", X"00", X"00", X"01", X"0f", X"00", X"08", X"00", X"41", X"2f", X"14", X"10", X"26", X"2f", X"43", X"2f", X"2b", X"28", X"26", X"00", X"0a", X"00", X"0b", X"12", X"22", X"02", X"02", X"03", X"09", X"05", X"00", X"03", X"16", X"12", X"26", X"19", X"32", X"0c", X"09", X"1c", X"25", X"20", X"25", X"20", X"29", X"3c", X"59", X"55", X"7f", X"7b", X"6f", X"4f", X"21", X"3a", X"2b", X"21", X"1b", X"00", X"2d", X"06", X"09", X"06", X"00", X"00", X"07", X"03", X"05", X"09", X"0a", X"05", X"04", X"00", X"39", X"2c", X"28", X"27", X"30", X"1d", X"33", X"2a", X"2c", X"3b", X"2f", X"00", X"1f", X"00", X"00", X"18", X"0a", X"05", X"03", X"19", X"0b", X"12", X"2a", X"0d", X"19", X"18", X"32", X"28", X"2d", X"2f", X"1e", X"02", X"00", X"1d", X"24", X"31", X"36", X"40", X"51", X"4e", X"6b", X"66", X"5b", X"3c", X"43", X"34", X"2d", X"24", X"1c", X"00", X"23", X"14", X"07", X"00", X"00", X"00", X"00", X"04", X"04", X"0a", X"13", X"00", X"06", X"02", X"6d", X"66", X"35", X"1e", X"10", X"1b", X"1a", X"3e", X"3f", X"4e", X"2d", X"18", X"14", X"00", X"1e", X"08", X"10", X"00", X"00", X"0b", X"0e", X"0e", X"2f", X"3c", X"4b", X"35", X"34", X"36", X"40", X"22", X"18", X"1a", X"0e", X"26", X"2f", X"34", X"26", X"43", X"3c", X"44", X"47", X"40", X"40", X"3d", X"4a", X"3b", X"2f", X"28", X"25", X"15", X"00", X"22", X"0a", X"02", X"05", X"05", X"00", X"00", X"03", X"03", X"0b", X"0e", X"01", X"00", X"68", X"4f", X"2c", X"22", X"34", X"25", X"27", X"37", X"45", X"30", X"43", X"3b", X"2a", X"4a", X"03", X"07", X"08", X"22", X"00", X"17", X"28", X"2a", X"24", X"31", X"28", X"38", X"2b", X"1c", X"28", X"26", X"32", X"29", X"26", X"2e", X"32", X"37", X"32", X"2e", X"45", X"6c", X"63", X"68", X"53", X"42", X"27", X"3e", X"3b", X"35", X"45", X"2a", X"15", X"00", X"1b", X"03", X"01", X"02", X"06", X"0d", X"03", X"00", X"0d", X"05", X"06", X"00", X"57", X"49", X"38", X"1c", X"47", X"20", X"2e", X"1c", X"1f", X"2b", X"30", X"38", X"27", X"2b", X"1a", X"07", X"10", X"17", X"06", X"1e", X"2b", X"27", X"28", X"22", X"31", X"32", X"35", X"3e", X"2f", X"2c", X"42", X"60", X"47", X"54", X"38", X"3d", X"39", X"1f", X"57", X"4f", X"6f", X"6c", X"3e", X"50", X"3e", X"35", X"3d", X"5d", X"39", X"30", X"2c", X"25", X"20", X"19", X"14", X"1a", X"2f", X"05", X"14", X"04", X"06", X"00", X"00", X"0f", X"6d", X"5e", X"51", X"45", X"38", X"36", X"33", X"48", X"25", X"32", X"34", X"4b", X"44", X"45", X"1f", X"05", X"2c", X"03", X"31", X"00", X"28", X"31", X"4c", X"31", X"56", X"76", X"61", X"72", X"4e", X"4d", X"51", X"39", X"4f", X"44", X"40", X"44", X"2d", X"13", X"26", X"4e", X"56", X"50", X"39", X"69", X"67", X"42", X"70", X"52", X"60", X"3c", X"39", X"33", X"35", X"41", X"2f", X"04", X"15", X"05", X"01", X"03", X"06", X"00", X"0c", X"06", X"6b", X"5a", X"4a", X"3c", X"16", X"1b", X"35", X"3f", X"31", X"58", X"4f", X"41", X"4f", X"38", X"3e", X"53", X"3a", X"41", X"37", X"36", X"3c", X"3f", X"3a", X"26", X"33", X"51", X"57", X"43", X"3e", X"5a", X"36", X"30", X"33", X"2d", X"2c", X"18", X"29", X"44", X"36", X"66", X"5d", X"5f", X"5a", X"53", X"5a", X"70", X"7e", X"64", X"36", X"49", X"40", X"3a", X"2e", X"0e", X"27", X"0d", X"03", X"02", X"07", X"00", X"00", X"08", X"05", X"02", X"7d", X"3e", X"62", X"40", X"2a", X"37", X"3f", X"2c", X"36", X"2d", X"2a", X"1f", X"3c", X"23", X"47", X"3d", X"46", X"5a", X"57", X"6e", X"49", X"3b", X"3f", X"13", X"31", X"25", X"2c", X"0f", X"46", X"3d", X"32", X"3b", X"23", X"3d", X"2b", X"23", X"25", X"1e", X"26", X"32", X"4c", X"3e", X"52", X"60", X"60", X"50", X"48", X"66", X"29", X"4a", X"43", X"34", X"15", X"2e", X"14", X"01", X"01", X"00", X"02", X"00", X"0e", X"05", X"01", X"00", X"7f", X"51", X"5f", X"5e", X"60", X"40", X"4a", X"32", X"36", X"0f", X"0f", X"1a", X"36", X"28", X"27", X"32", X"3c", X"43", X"59", X"5d", X"32", X"36", X"3d", X"1e", X"13", X"20", X"0a", X"0f", X"2c", X"26", X"32", X"47", X"30", X"3e", X"45", X"1e", X"25", X"0d", X"18", X"39", X"31", X"4b", X"50", X"41", X"44", X"58", X"51", X"71", X"54", X"5b", X"3f", X"26", X"00", X"24", X"0d", X"03", X"04", X"03", X"05", X"00", X"05", X"03", X"00", X"00", X"55", X"47", X"68", X"44", X"37", X"2b", X"39", X"18", X"29", X"00", X"00", X"1c", X"3e", X"1e", X"27", X"25", X"3b", X"3d", X"2a", X"2a", X"34", X"32", X"3d", X"27", X"0e", X"12", X"00", X"01", X"00", X"02", X"29", X"29", X"54", X"33", X"2f", X"2a", X"20", X"11", X"07", X"1b", X"29", X"2c", X"27", X"1e", X"25", X"36", X"3c", X"52", X"4f", X"48", X"45", X"22", X"00", X"29", X"0e", X"00", X"01", X"01", X"04", X"00", X"03", X"00", X"01", X"00", X"44", X"2a", X"54", X"42", X"40", X"34", X"30", X"30", X"1e", X"05", X"17", X"23", X"2e", X"29", X"38", X"3b", X"51", X"51", X"31", X"3c", X"35", X"55", X"2e", X"16", X"17", X"00", X"00", X"17", X"09", X"04", X"17", X"1b", X"2f", X"32", X"34", X"35", X"23", X"2c", X"07", X"05", X"05", X"16", X"2c", X"16", X"31", X"30", X"28", X"21", X"32", X"37", X"4b", X"3a", X"26", X"00", X"16", X"03", X"00", X"03", X"00", X"00", X"07", X"00", X"00", X"02", X"3f", X"52", X"47", X"44", X"39", X"3a", X"21", X"21", X"24", X"33", X"4b", X"2b", X"18", X"1b", X"25", X"23", X"23", X"21", X"2a", X"25", X"1c", X"1b", X"13", X"00", X"11", X"05", X"01", X"16", X"17", X"04", X"05", X"07", X"24", X"39", X"32", X"37", X"2c", X"3c", X"03", X"07", X"06", X"1a", X"2a", X"24", X"24", X"3a", X"31", X"42", X"46", X"3d", X"54", X"47", X"40", X"29", X"00", X"23", X"10", X"00", X"04", X"00", X"00", X"0a", X"06", X"04", X"46", X"4a", X"52", X"78", X"4b", X"51", X"41", X"53", X"70", X"47", X"4e", X"65", X"37", X"29", X"41", X"1f", X"25", X"00", X"03", X"16", X"1e", X"10", X"03", X"12", X"0a", X"00", X"07", X"06", X"0f", X"08", X"00", X"33", X"33", X"0f", X"2f", X"3d", X"3a", X"33", X"03", X"0c", X"10", X"16", X"2c", X"1f", X"2f", X"06", X"1e", X"2f", X"41", X"3e", X"44", X"34", X"32", X"29", X"29", X"2d", X"00", X"19", X"0c", X"02", X"00", X"0c", X"03", X"00", X"4d", X"50", X"4e", X"4e", X"68", X"48", X"4c", X"67", X"5f", X"4a", X"6b", X"58", X"38", X"37", X"35", X"12", X"18", X"1e", X"23", X"2c", X"23", X"18", X"30", X"2a", X"1e", X"25", X"24", X"0a", X"0f", X"0f", X"01", X"0f", X"16", X"21", X"2d", X"44", X"69", X"2a", X"27", X"19", X"22", X"1a", X"34", X"3f", X"3c", X"2c", X"4e", X"55", X"65", X"70", X"56", X"35", X"15", X"29", X"24", X"12", X"1c", X"00", X"07", X"15", X"0d", X"00", X"08", X"01", X"33", X"31", X"33", X"44", X"4a", X"78", X"7c", X"46", X"5e", X"7b", X"42", X"5e", X"68", X"76", X"5a", X"62", X"44", X"4f", X"34", X"37", X"2e", X"35", X"3c", X"33", X"2d", X"2e", X"32", X"19", X"1c", X"06", X"06", X"0c", X"3e", X"14", X"2a", X"2f", X"3b", X"4a", X"4d", X"50", X"4e", X"44", X"4b", X"37", X"42", X"50", X"3d", X"65", X"56", X"43", X"45", X"10", X"31", X"13", X"0a", X"07", X"07", X"06", X"11", X"00", X"06", X"01", X"00", X"0f", X"1b", X"23", X"28", X"37", X"41", X"65", X"56", X"3d", X"54", X"61", X"40", X"59", X"68", X"5a", X"51", X"69", X"43", X"44", X"4d", X"6d", X"5f", X"44", X"30", X"24", X"23", X"29", X"2c", X"26", X"10", X"05", X"08", X"01", X"0c", X"1c", X"3a", X"32", X"34", X"23", X"22", X"31", X"33", X"30", X"34", X"44", X"28", X"3f", X"61", X"4c", X"3e", X"37", X"23", X"00", X"21", X"0f", X"07", X"02", X"01", X"01", X"00", X"03", X"11", X"12", X"10", X"00", X"0c", X"13", X"25", X"34", X"58", X"32", X"49", X"20", X"3d", X"5f", X"4f", X"54", X"4a", X"4f", X"60", X"6b", X"76", X"6b", X"71", X"69", X"60", X"4b", X"54", X"4e", X"49", X"29", X"2e", X"36", X"38", X"15", X"09", X"00", X"12", X"0d", X"2b", X"31", X"2c", X"2c", X"2e", X"38", X"39", X"32", X"34", X"09", X"3b", X"52", X"52", X"50", X"3d", X"35", X"2a", X"01", X"18", X"08", X"05", X"01", X"00", X"00", X"00", X"04", X"04", X"03", X"03", X"0f", X"32", X"00", X"17", X"2a", X"38", X"3c", X"3f", X"4d", X"35", X"3a", X"74", X"7f", X"7e", X"40", X"57", X"69", X"6c", X"5e", X"69", X"6c", X"52", X"4a", X"4a", X"4f", X"51", X"3e", X"4d", X"4c", X"4d", X"35", X"17", X"03", X"00", X"13", X"1f", X"2c", X"2b", X"3a", X"37", X"31", X"39", X"45", X"3a", X"1e", X"3a", X"56", X"74", X"7b", X"71", X"5b", X"41", X"37", X"00", X"20", X"0a", X"01", X"04", X"09", X"01", X"10", X"02", X"00", X"00", X"09", X"32", X"00", X"1c", X"3a", X"41", X"41", X"41", X"46", X"30", X"61", X"74", X"70", X"7b", X"7c", X"64", X"6d", X"5e", X"56", X"53", X"5f", X"4f", X"4e", X"39", X"3d", X"3c", X"42", X"47", X"4a", X"3b", X"1e", X"1d", X"12", X"12", X"10", X"29", X"10", X"21", X"3a", X"28", X"3b", X"3d", X"32", X"38", X"2e", X"38", X"50", X"58", X"4a", X"4f", X"38", X"3a", X"2b", X"2b", X"27", X"2f", X"36", X"07", X"14", X"0b", X"00", X"08", X"01", X"02", X"02", X"29", X"00", X"21", X"3b", X"3e", X"3a", X"3a", X"35", X"5b", X"6b", X"64", X"75", X"69", X"50", X"5e", X"58", X"4c", X"4c", X"76", X"58", X"5d", X"5c", X"51", X"43", X"4f", X"3d", X"43", X"2f", X"1f", X"0a", X"04", X"06", X"08", X"15", X"16", X"24", X"0e", X"29", X"38", X"67", X"36", X"26", X"4a", X"2c", X"3e", X"3a", X"5d", X"4f", X"20", X"49", X"44", X"41", X"37", X"17", X"1b", X"13", X"0a", X"00", X"00", X"0a", X"00", X"00", X"03", X"02", X"3b", X"13", X"34", X"38", X"35", X"38", X"3c", X"4d", X"33", X"3f", X"72", X"6b", X"69", X"4f", X"55", X"61", X"65", X"30", X"45", X"55", X"5e", X"5f", X"5a", X"44", X"42", X"3a", X"52", X"35", X"2e", X"2f", X"28", X"27", X"09", X"1b", X"15", X"1f", X"21", X"3e", X"2b", X"2d", X"25", X"19", X"0f", X"24", X"52", X"61", X"40", X"57", X"25", X"45", X"3a", X"36", X"33", X"25", X"01", X"1a", X"0a", X"00", X"06", X"02", X"00", X"01", X"03", X"00", X"19", X"3e", X"2a", X"21", X"22", X"22", X"1e", X"2a", X"32", X"64", X"46", X"3c", X"37", X"49", X"4a", X"51", X"56", X"5f", X"3f", X"51", X"60", X"62", X"56", X"52", X"5d", X"66", X"72", X"71", X"2d", X"28", X"29", X"13", X"11", X"0c", X"05", X"3b", X"38", X"34", X"14", X"2e", X"10", X"25", X"3c", X"48", X"47", X"37", X"7f", X"75", X"57", X"38", X"45", X"33", X"2e", X"24", X"0e", X"1a", X"10", X"1a", X"0d", X"03", X"01", X"00", X"00", X"00", X"27", X"04", X"1d", X"0d", X"0a", X"15", X"27", X"32", X"52", X"33", X"3f", X"41", X"1d", X"2c", X"39", X"47", X"52", X"64", X"3a", X"4e", X"58", X"58", X"57", X"62", X"6c", X"74", X"78", X"6b", X"20", X"1b", X"0f", X"00", X"0a", X"10", X"21", X"0c", X"23", X"3a", X"29", X"28", X"1c", X"1a", X"5a", X"4e", X"49", X"7e", X"76", X"68", X"5c", X"41", X"36", X"27", X"1b", X"2e", X"14", X"03", X"01", X"00", X"0e", X"00", X"07", X"00", X"00", X"00", X"01", X"03", X"02", X"10", X"22", X"00", X"11", X"22", X"25", X"2b", X"30", X"2d", X"3d", X"19", X"31", X"3f", X"4e", X"57", X"3e", X"4d", X"61", X"66", X"6b", X"5f", X"73", X"75", X"71", X"42", X"29", X"1f", X"15", X"0b", X"00", X"1b", X"20", X"23", X"2c", X"37", X"18", X"32", X"35", X"43", X"5c", X"5f", X"53", X"44", X"4c", X"3e", X"22", X"3d", X"2b", X"14", X"00", X"15", X"09", X"00", X"00", X"00", X"04", X"05", X"01", X"03", X"00", X"00", X"01", X"03", X"04", X"02", X"06", X"18", X"00", X"15", X"24", X"29", X"33", X"39", X"41", X"3d", X"34", X"4b", X"3f", X"4d", X"65", X"70", X"76", X"74", X"5d", X"52", X"56", X"48", X"42", X"3d", X"49", X"3b", X"0f", X"1c", X"0d", X"15", X"1c", X"20", X"2e", X"45", X"2a", X"20", X"2b", X"58", X"55", X"64", X"72", X"69", X"4b", X"43", X"3d", X"3d", X"2c", X"15", X"00", X"28", X"0a", X"00", X"04", X"02", X"08", X"08", X"02", X"00", X"04", X"02", X"01", X"03", X"04", X"03", X"06", X"19", X"00", X"1b", X"22", X"2a", X"2d", X"34", X"3a", X"3a", X"38", X"4a", X"4e", X"62", X"6d", X"73", X"72", X"70", X"6d", X"59", X"55", X"55", X"56", X"38", X"3a", X"35", X"1e", X"05", X"12", X"3f", X"3f", X"2f", X"38", X"1c", X"0c", X"26", X"3b", X"3e", X"57", X"48", X"6d", X"67", X"42", X"4b", X"23", X"40", X"39", X"27", X"1d", X"00", X"1a", X"08", X"11", X"00", X"09", X"00", X"0a", X"06", X"04", X"05", X"00", X"04", X"01", X"06", X"0a", X"1d", X"01", X"1b", X"1f", X"27", X"2c", X"38", X"3b", X"19", X"35", X"47", X"62", X"47", X"62", X"71", X"78", X"7b", X"72", X"6d", X"53", X"55", X"5c", X"34", X"31", X"17", X"0b", X"15", X"28", X"3a", X"2e", X"1b", X"1d", X"03", X"0f", X"15", X"2d", X"54", X"6b", X"7b", X"58", X"4a", X"58", X"58", X"4c", X"3f", X"59", X"46", X"30", X"2b", X"2a", X"31", X"00", X"1c", X"0b", X"02", X"01", X"02", X"0a", X"16", X"02", X"05", X"03", X"07", X"17", X"00", X"1d", X"26", X"29", X"2f", X"34", X"3d", X"19", X"39", X"45", X"5a", X"5e", X"64", X"69", X"6c", X"6f", X"6c", X"68", X"50", X"56", X"56", X"56", X"2d", X"21", X"21", X"43", X"1a", X"2d", X"20", X"20", X"31", X"17", X"0e", X"0d", X"1c", X"26", X"58", X"64", X"56", X"64", X"5a", X"52", X"3f", X"56", X"78", X"66", X"43", X"45", X"3e", X"38", X"00", X"1a", X"04", X"03", X"0b", X"07", X"03", X"00", X"04", X"06", X"11", X"1d", X"08", X"06", X"19", X"2a", X"35", X"58", X"4b", X"43", X"44", X"40", X"54", X"5a", X"5b", X"62", X"6c", X"41", X"51", X"53", X"4f", X"53", X"56", X"45", X"47", X"48", X"44", X"36", X"13", X"30", X"2f", X"34", X"32", X"1e", X"56", X"1d", X"09", X"10", X"2a", X"24", X"2d", X"37", X"47", X"48", X"53", X"58", X"60", X"56", X"7f", X"55", X"33", X"4e", X"34", X"0c", X"33", X"13", X"09", X"04", X"02", X"00", X"08", X"01", X"00", X"14", X"07", X"2f", X"41", X"3a", X"37", X"35", X"37", X"3a", X"34", X"59", X"77", X"71", X"70", X"6a", X"6e", X"71", X"74", X"75", X"3c", X"47", X"56", X"66", X"75", X"79", X"6e", X"58", X"2f", X"27", X"0f", X"12", X"17", X"34", X"32", X"4a", X"46", X"12", X"07", X"1c", X"09", X"17", X"2d", X"3c", X"3b", X"4c", X"56", X"70", X"50", X"58", X"5e", X"49", X"5f", X"4c", X"38", X"18", X"1f", X"16", X"07", X"09", X"04", X"0c", X"11", X"06", X"00", X"01", X"09", X"09", X"1b", X"0e", X"2e", X"3a", X"3e", X"3e", X"41", X"37", X"44", X"59", X"7b", X"7c", X"79", X"72", X"63", X"7f", X"40", X"50", X"52", X"48", X"55", X"71", X"77", X"60", X"31", X"1e", X"1a", X"26", X"27", X"3e", X"31", X"34", X"4c", X"37", X"09", X"04", X"11", X"18", X"39", X"3e", X"31", X"2f", X"3e", X"34", X"2d", X"48", X"3f", X"55", X"55", X"3e", X"45", X"41", X"2a", X"05", X"1f", X"13", X"06", X"00", X"00", X"03", X"0a", X"00", X"0c", X"11", X"01", X"22", X"30", X"34", X"38", X"3b", X"40", X"4c", X"27", X"56", X"44", X"75", X"75", X"7e", X"7e", X"48", X"42", X"4b", X"53", X"45", X"4f", X"4d", X"43", X"27", X"29", X"2a", X"10", X"19", X"07", X"23", X"2e", X"32", X"20", X"28", X"21", X"06", X"07", X"0c", X"0c", X"26", X"23", X"1d", X"0c", X"17", X"29", X"1f", X"35", X"23", X"3d", X"3e", X"36", X"4e", X"33", X"00", X"28", X"17", X"00", X"08", X"05", X"01", X"00", X"27", X"10", X"16", X"21", X"2b", X"33", X"38", X"3b", X"3f", X"42", X"49", X"22", X"47", X"5f", X"55", X"4d", X"59", X"3a", X"40", X"4a", X"55", X"50", X"3e", X"49", X"45", X"3d", X"3c", X"22", X"0c", X"0b", X"0a", X"2f", X"59", X"3e", X"21", X"2a", X"2f", X"41", X"2b", X"04", X"00", X"0a", X"0f", X"11", X"05", X"30", X"2c", X"38", X"3a", X"39", X"30", X"27", X"35", X"36", X"3a", X"1e", X"23", X"09", X"05", X"09", X"10", X"04", X"03", X"02", X"03", X"04", X"01", X"14", X"00", X"1c", X"2c", X"34", X"39", X"3f", X"49", X"2c", X"42", X"5d", X"44", X"61", X"51", X"69", X"50", X"60", X"4d", X"3f", X"47", X"4b", X"41", X"49", X"44", X"20", X"15", X"18", X"2a", X"36", X"44", X"3b", X"22", X"37", X"4b", X"55", X"43", X"21", X"17", X"00", X"00", X"16", X"0d", X"13", X"1f", X"2f", X"4a", X"35", X"3f", X"42", X"4c", X"2c", X"52", X"27", X"27", X"21", X"05", X"00", X"05", X"00", X"03", X"00", X"02", X"02", X"00", X"10", X"15", X"0a", X"40", X"40", X"2b", X"2b", X"39", X"49", X"56", X"64", X"63", X"5d", X"6c", X"66", X"56", X"63", X"71", X"54", X"5d", X"5a", X"50", X"23", X"11", X"06", X"18", X"24", X"3a", X"3b", X"4c", X"3e", X"37", X"31", X"14", X"28", X"2c", X"1e", X"20", X"0f", X"0e", X"12", X"2c", X"1d", X"13", X"2f", X"05", X"0e", X"2a", X"29", X"36", X"47", X"61", X"40", X"40", X"19", X"1e", X"00", X"08", X"08", X"00", X"00", X"00", X"00", X"07", X"14", X"2d", X"00", X"16", X"2d", X"60", X"6e", X"45", X"62", X"63", X"6f", X"3d", X"54", X"6b", X"6c", X"5a", X"66", X"75", X"72", X"40", X"41", X"2b", X"27", X"07", X"16", X"40", X"11", X"22", X"23", X"28", X"38", X"26", X"36", X"32", X"33", X"3e", X"48", X"40", X"50", X"47", X"38", X"46", X"3c", X"24", X"1e", X"15", X"10", X"37", X"26", X"22", X"42", X"44", X"3e", X"44", X"09", X"21", X"0c", X"0d", X"00", X"04", X"02", X"00", X"02", X"00", X"13", X"14", X"06", X"1b", X"34", X"42", X"72", X"78", X"60", X"60", X"56", X"5c", X"59", X"6c", X"3d", X"44", X"4d", X"69", X"4f", X"4b", X"30", X"1d", X"07", X"00", X"20", X"42", X"1f", X"3d", X"4f", X"3f", X"39", X"2b", X"38", X"30", X"48", X"2b", X"1d", X"27", X"3c", X"2f", X"2d", X"28", X"33", X"31", X"29", X"45", X"34", X"2b", X"1b", X"2d", X"1a", X"22", X"35", X"35", X"1e", X"2a", X"04", X"07", X"00", X"00", X"00", X"22", X"0a", X"09", X"0a", X"19", X"2c", X"2e", X"36", X"45", X"5c", X"7a", X"7f", X"60", X"6d", X"6b", X"51", X"45", X"49", X"3f", X"3d", X"35", X"31", X"36", X"38", X"0c", X"12", X"02", X"10", X"2a", X"2d", X"39", X"43", X"65", X"74", X"3c", X"4e", X"27", X"39", X"08", X"0d", X"0e", X"22", X"2e", X"2a", X"34", X"1c", X"5d", X"53", X"4c", X"61", X"34", X"2f", X"42", X"2b", X"19", X"2a", X"34", X"27", X"22", X"00", X"03", X"05", X"01", X"00", X"21", X"00", X"35", X"3c", X"3f", X"3d", X"43", X"4c", X"4b", X"55", X"65", X"40", X"5a", X"64", X"4a", X"58", X"2f", X"2a", X"17", X"2b", X"26", X"16", X"17", X"00", X"00", X"0c", X"03", X"32", X"28", X"35", X"3a", X"33", X"19", X"1a", X"4e", X"3a", X"30", X"45", X"1f", X"03", X"00", X"0c", X"20", X"28", X"31", X"5e", X"4b", X"62", X"78", X"4f", X"47", X"49", X"4a", X"47", X"61", X"59", X"33", X"19", X"1d", X"05", X"02", X"01", X"06", X"02", X"00", X"18", X"13", X"4a", X"41", X"4d", X"5c", X"75", X"4f", X"62", X"66", X"55", X"68", X"6b", X"53", X"2f", X"2b", X"20", X"2c", X"08", X"09", X"03", X"13", X"1a", X"19", X"19", X"34", X"3d", X"3d", X"34", X"26", X"24", X"04", X"22", X"28", X"28", X"22", X"2a", X"15", X"1e", X"33", X"51", X"51", X"46", X"4d", X"4e", X"7f", X"4f", X"41", X"63", X"56", X"42", X"4c", X"58", X"34", X"1b", X"0f", X"24", X"15", X"00", X"00", X"00", X"00", X"00", X"04", X"1e", X"10", X"38", X"50", X"51", X"63", X"5b", X"53", X"5b", X"6b", X"4a", X"4d", X"5b", X"35", X"2d", X"3f", X"21", X"1c", X"2c", X"1f", X"24", X"20", X"20", X"25", X"2e", X"2f", X"34", X"3d", X"21", X"3c", X"0a", X"00", X"0f", X"22", X"36", X"2e", X"42", X"31", X"13", X"3e", X"4e", X"60", X"4b", X"7e", X"54", X"47", X"3c", X"34", X"2e", X"2d", X"46", X"2c", X"2b", X"0d", X"19", X"0a", X"06", X"12", X"0d", X"00", X"00", X"02", X"00", X"2f", X"0a", X"32", X"42", X"35", X"38", X"34", X"2c", X"38", X"3d", X"3d", X"3c", X"30", X"3b", X"2e", X"26", X"38", X"3f", X"3c", X"24", X"39", X"29", X"25", X"42", X"31", X"3a", X"2d", X"35", X"28", X"1e", X"17", X"1c", X"20", X"2c", X"49", X"18", X"2d", X"3a", X"2a", X"4c", X"5d", X"47", X"64", X"49", X"59", X"3e", X"52", X"32", X"15", X"30", X"0a", X"2c", X"2d", X"20", X"04", X"01", X"0b", X"0d", X"0d", X"04", X"07", X"01", X"01", X"00", X"26", X"3f", X"45", X"2c", X"27", X"33", X"2e", X"1e", X"26", X"27", X"32", X"0f", X"09", X"17", X"2d", X"39", X"32", X"39", X"2f", X"50", X"23", X"07", X"04", X"0b", X"03", X"25", X"18", X"30", X"1d", X"1d", X"34", X"41", X"46", X"3f", X"2e", X"14", X"0e", X"27", X"31", X"42", X"5f", X"41", X"3e", X"42", X"3b", X"3a", X"39", X"26", X"1d", X"22", X"23", X"00", X"12", X"0b", X"0c", X"00", X"00", X"02", X"02", X"03", X"0e", X"05", X"02", X"00", X"33", X"00", X"38", X"58", X"39", X"47", X"3a", X"2d", X"35", X"31", X"26", X"3b", X"0e", X"42", X"32", X"3c", X"2c", X"4a", X"17", X"0a", X"03", X"14", X"20", X"1f", X"31", X"1c", X"2d", X"33", X"37", X"4b", X"5b", X"58", X"54", X"5f", X"4a", X"5e", X"35", X"2a", X"27", X"36", X"4c", X"7f", X"65", X"39", X"2a", X"2d", X"41", X"1e", X"00", X"14", X"10", X"07", X"09", X"03", X"18", X"00", X"00", X"03", X"01", X"06", X"04", X"00", X"02", X"00", X"33", X"00", X"27", X"47", X"48", X"42", X"3c", X"27", X"30", X"54", X"3c", X"41", X"28", X"10", X"22", X"2c", X"1d", X"11", X"0b", X"1f", X"2d", X"43", X"31", X"2b", X"40", X"45", X"3c", X"40", X"67", X"59", X"61", X"5b", X"53", X"68", X"69", X"4c", X"51", X"32", X"2c", X"33", X"37", X"43", X"4d", X"23", X"10", X"2b", X"00", X"25", X"02", X"0e", X"04", X"00", X"00", X"20", X"00", X"20", X"00", X"00", X"00", X"03", X"04", X"0e", X"04", X"00", X"0b", X"21", X"3a", X"2d", X"5b", X"3d", X"26", X"0f", X"2e", X"29", X"3c", X"3c", X"6c", X"74", X"39", X"36", X"2d", X"2a", X"14", X"1b", X"19", X"2d", X"3e", X"67", X"4f", X"39", X"44", X"57", X"54", X"67", X"64", X"43", X"7f", X"3e", X"54", X"7a", X"50", X"4a", X"57", X"49", X"68", X"52", X"46", X"01", X"18", X"0e", X"15", X"00", X"0a", X"00", X"0a", X"03", X"00", X"08", X"07", X"00", X"00", X"1e", X"01", X"02", X"00", X"0b", X"05", X"00", X"37", X"4c", X"58", X"54", X"5a", X"5a", X"35", X"18", X"28", X"0c", X"2b", X"3d", X"31", X"27", X"3a", X"2a", X"15", X"16", X"1f", X"23", X"4e", X"5f", X"4b", X"6a", X"70", X"64", X"6d", X"76", X"51", X"47", X"57", X"67", X"7f", X"6e", X"57", X"4c", X"4c", X"79", X"42", X"4c", X"3e", X"31", X"32", X"1f", X"1f", X"14", X"11", X"0a", X"04", X"08", X"02", X"03", X"07", X"00", X"31", X"00", X"00", X"01", X"00", X"0f", X"14", X"06", X"0d", X"00", X"2b", X"46", X"41", X"3b", X"3d", X"39", X"0e", X"20", X"2d", X"34", X"2d", X"32", X"33", X"2d", X"30", X"36", X"24", X"12", X"3d", X"47", X"59", X"4f", X"46", X"55", X"47", X"5a", X"65", X"64", X"50", X"67", X"65", X"40", X"71", X"5e", X"2b", X"36", X"2f", X"2f", X"35", X"3f", X"25", X"01", X"37", X"00", X"00", X"19", X"11", X"02", X"00", X"02", X"00", X"00", X"00", X"04", X"01", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"03", X"32", X"53", X"4b", X"45", X"41", X"23", X"2a", X"3a", X"48", X"3b", X"39", X"1d", X"46", X"33", X"2b", X"1e", X"1f", X"0d", X"2a", X"3f", X"4a", X"42", X"53", X"4e", X"6a", X"46", X"4e", X"5c", X"6b", X"5a", X"4d", X"4a", X"54", X"57", X"36", X"26", X"1f", X"1a", X"2d", X"30", X"04", X"22", X"0f", X"04", X"08", X"00", X"10", X"21", X"0b", X"00", X"00", X"00", X"00", X"00", X"00", X"2d", X"0d", X"10", X"0f", X"10", X"0f", X"00", X"00", X"0e", X"37", X"36", X"40", X"44", X"46", X"28", X"39", X"42", X"4c", X"38", X"49", X"37", X"3b", X"1e", X"1d", X"40", X"1c", X"2a", X"2c", X"5d", X"4f", X"4a", X"57", X"50", X"38", X"7f", X"7c", X"7a", X"3d", X"54", X"30", X"4d", X"4b", X"2b", X"2e", X"1f", X"04", X"47", X"49", X"00", X"0c", X"23", X"09", X"01", X"00", X"00", X"00", X"07", X"1b", X"00", X"00", X"04", X"03", X"00", X"0b", X"0d", X"0e", X"10", X"11", X"0d", X"11", X"0d", X"08", X"05", X"75", X"6c", X"51", X"49", X"40", X"3a", X"23", X"00", X"0d", X"0a", X"0a", X"2b", X"1d", X"2b", X"2c", X"2b", X"1d", X"1c", X"2f", X"69", X"74", X"62", X"49", X"43", X"64", X"66", X"77", X"78", X"75", X"4b", X"24", X"42", X"3c", X"33", X"29", X"14", X"26", X"06", X"11", X"17", X"00", X"24", X"0c", X"00", X"00", X"0e", X"0b", X"03", X"00", X"1d", X"05", X"04", X"00", X"00", X"0a", X"0c", X"0b", X"08", X"11", X"10", X"11", X"10", X"0f", X"0e", X"58", X"4b", X"43", X"28", X"27", X"27", X"1a", X"00", X"01", X"12", X"00", X"1e", X"34", X"4c", X"2d", X"32", X"2e", X"2f", X"38", X"3e", X"4f", X"46", X"53", X"4d", X"38", X"77", X"6e", X"6f", X"74", X"53", X"33", X"43", X"3e", X"42", X"33", X"06", X"17", X"03", X"01", X"09", X"0f", X"0c", X"04", X"00", X"06", X"00", X"03", X"03", X"00", X"00", X"00", X"2d", X"00", X"0f", X"0e", X"0f", X"0f", X"12", X"0c", X"0e", X"10", X"0f", X"0c", X"0a"
    );

begin

    process(video_on, R_int, G_int, B_int)
    begin
        if (video_on = '1') then
            R <= R_int(6 downto 0);
            G <= G_int(6 downto 0);
            B <= B_int(6 downto 0);
        else
            R <= (others => '0');
            G <= (others => '0');
            B <= (others => '0');
        end if;
    end process;

    -- ROM
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (re = '1') then
                R_int <= r_rom(to_integer(unsigned(pixel_y) * 64 + unsigned(pixel_x)));
                G_int <= g_rom(to_integer(unsigned(pixel_y) * 64 + unsigned(pixel_x)));
                B_int <= b_rom(to_integer(unsigned(pixel_y) * 64 + unsigned(pixel_x)));
            end if;
        end if;
    end process;

end Behavioral;

